module Signed(output [31:0] AnswerOne,output [31:0] AnswerTwo,input [31:0] A,input [31:0] B,input OpCode);

endmodule