//Define 32 bit multiplexer
module UMultiplier(O, X, Y);

// I/O port declaration
input [31:0] X, Y;
output [63:0] O;

//internal nets

wire [1023:0] C;
wire [639:0]sum, carry; 
wire [447:0] sum_1,carry_1;
wire [319:0] sum_2,carry_2;
wire [191:0] sum_3,carry_3;
wire [127:0] sum_4,carry_4;
wire [63:0] sum_5,carry_5;
wire [63:0] sum_6,carry_6;
wire [63:0] sum_7,carry_7;
wire [63:0] carry_8;

//Instantiate logic gate primitives

//1.1

//PP0
and (C[0], X[0], Y[0]);
and (C[1], X[1], Y[0]);
and (C[2], X[2], Y[0]);
and (C[3], X[3], Y[0]);
and (C[4], X[4], Y[0]);
and (C[5], X[5], Y[0]);
and (C[6], X[6], Y[0]);
and (C[7], X[7], Y[0]);
and (C[8], X[8], Y[0]);
and (C[9], X[9], Y[0]);
and (C[10], X[10], Y[0]);
and (C[11], X[11], Y[0]);
and (C[12], X[12], Y[0]);
and (C[13], X[13], Y[0]);
and (C[14], X[14], Y[0]);
and (C[15], X[15], Y[0]);
and (C[16], X[16], Y[0]);
and (C[17], X[17], Y[0]);
and (C[18], X[18], Y[0]);
and (C[19], X[19], Y[0]);
and (C[20], X[20], Y[0]);
and (C[21], X[21], Y[0]);
and (C[22], X[22], Y[0]);
and (C[23], X[23], Y[0]);
and (C[24], X[24], Y[0]);
and (C[25], X[25], Y[0]);
and (C[26], X[26], Y[0]);
and (C[27], X[27], Y[0]);
and (C[28], X[28], Y[0]);
and (C[29], X[29], Y[0]);
and (C[30], X[30], Y[0]);
and (C[31], X[31], Y[0]);

//PP1

and (C[32], X[0], Y[1]);
and (C[33], X[1], Y[1]);
and (C[34], X[2], Y[1]);
and (C[35], X[3], Y[1]);
and (C[36], X[4], Y[1]);
and (C[37], X[5], Y[1]);
and (C[38], X[6], Y[1]);
and (C[39], X[7], Y[1]);
and (C[40], X[8], Y[1]);
and (C[41], X[9], Y[1]);
and (C[42], X[10], Y[1]);
and (C[43], X[11], Y[1]);
and (C[44], X[12], Y[1]);
and (C[45], X[13], Y[1]);
and (C[46], X[14], Y[1]);
and (C[47], X[15], Y[1]);
and (C[48], X[16], Y[1]);
and (C[49], X[17], Y[1]);
and (C[50], X[18], Y[1]);
and (C[51], X[19], Y[1]);
and (C[52], X[20], Y[1]);
and (C[53], X[21], Y[1]);
and (C[54], X[22], Y[1]);
and (C[55], X[23], Y[1]);
and (C[56], X[24], Y[1]);
and (C[57], X[25], Y[1]);
and (C[58], X[26], Y[1]);
and (C[59], X[27], Y[1]);
and (C[60], X[28], Y[1]);
and (C[61], X[29], Y[1]);
and (C[62], X[30], Y[1]);
and (C[63], X[31], Y[1]);

//PP2
and (C[64], X[0], Y[2]);
and (C[65], X[1], Y[2]);
and (C[66], X[2], Y[2]);
and (C[67], X[3], Y[2]);
and (C[68], X[4], Y[2]);
and (C[69], X[5], Y[2]);
and (C[70], X[6], Y[2]);
and (C[71], X[7], Y[2]);
and (C[72], X[8], Y[2]);
and (C[73], X[9], Y[2]);
and (C[74], X[10], Y[2]);
and (C[75], X[11], Y[2]);
and (C[76], X[12], Y[2]);
and (C[77], X[13], Y[2]);
and (C[78], X[14], Y[2]);
and (C[79], X[15], Y[2]);
and (C[80], X[16], Y[2]);
and (C[81], X[17], Y[2]);
and (C[82], X[18], Y[2]);
and (C[83], X[19], Y[2]);
and (C[84], X[20], Y[2]);
and (C[85], X[21], Y[2]);
and (C[86], X[22], Y[2]);
and (C[87], X[23], Y[2]);
and (C[88], X[24], Y[2]);
and (C[89], X[25], Y[2]);
and (C[90], X[26], Y[2]);
and (C[91], X[27], Y[2]);
and (C[92], X[28], Y[2]);
and (C[93], X[29], Y[2]);
and (C[94], X[30], Y[2]);
and (C[95], X[31], Y[2]);

//PP3
and (C[96], X[0], Y[3]);
and (C[97], X[1], Y[3]);
and (C[98], X[2], Y[3]);
and (C[99], X[3], Y[3]);
and (C[100], X[4], Y[3]);
and (C[101], X[5], Y[3]);
and (C[102], X[6], Y[3]);
and (C[103], X[7], Y[3]);
and (C[104], X[8], Y[3]);
and (C[105], X[9], Y[3]);
and (C[106], X[10], Y[3]);
and (C[107], X[11], Y[3]);
and (C[108], X[12], Y[3]);
and (C[109], X[13], Y[3]);
and (C[110], X[14], Y[3]);
and (C[111], X[15], Y[3]);
and (C[112], X[16], Y[3]);
and (C[113], X[17], Y[3]);
and (C[114], X[18], Y[3]);
and (C[115], X[19], Y[3]);
and (C[116], X[20], Y[3]);
and (C[117], X[21], Y[3]);
and (C[118], X[22], Y[3]);
and (C[119], X[23], Y[3]);
and (C[120], X[24], Y[3]);
and (C[121], X[25], Y[3]);
and (C[122], X[26], Y[3]);
and (C[123], X[27], Y[3]);
and (C[124], X[28], Y[3]);
and (C[125], X[29], Y[3]);
and (C[126], X[30], Y[3]);
and (C[127], X[31], Y[3]);

//PP4
and (C[128], X[0], Y[4]);
and (C[129], X[1], Y[4]);
and (C[130], X[2], Y[4]);
and (C[131], X[3], Y[4]);
and (C[132], X[4], Y[4]);
and (C[133], X[5], Y[4]);
and (C[134], X[6], Y[4]);
and (C[135], X[7], Y[4]);
and (C[136], X[8], Y[4]);
and (C[137], X[9], Y[4]);
and (C[138], X[10], Y[4]);
and (C[139], X[11], Y[4]);
and (C[140], X[12], Y[4]);
and (C[141], X[13], Y[4]);
and (C[142], X[14], Y[4]);
and (C[143], X[15], Y[4]);
and (C[144], X[16], Y[4]);
and (C[145], X[17], Y[4]);
and (C[146], X[18], Y[4]);
and (C[147], X[19], Y[4]);
and (C[148], X[20], Y[4]);
and (C[149], X[21], Y[4]);
and (C[150], X[22], Y[4]);
and (C[151], X[23], Y[4]);
and (C[152], X[24], Y[4]);
and (C[153], X[25], Y[4]);
and (C[154], X[26], Y[4]);
and (C[155], X[27], Y[4]);
and (C[156], X[28], Y[4]);
and (C[157], X[29], Y[4]);
and (C[158], X[30], Y[4]);
and (C[159], X[31], Y[4]);

//PP5
and (C[160], X[0], Y[5]);
and (C[161], X[1], Y[5]);
and (C[162], X[2], Y[5]);
and (C[163], X[3], Y[5]);
and (C[164], X[4], Y[5]);
and (C[165], X[5], Y[5]);
and (C[166], X[6], Y[5]);
and (C[167], X[7], Y[5]);
and (C[168], X[8], Y[5]);
and (C[169], X[9], Y[5]);
and (C[170], X[10], Y[5]);
and (C[171], X[11], Y[5]);
and (C[172], X[12], Y[5]);
and (C[173], X[13], Y[5]);
and (C[174], X[14], Y[5]);
and (C[175], X[15], Y[5]);
and (C[176], X[16], Y[5]);
and (C[177], X[17], Y[5]);
and (C[178], X[18], Y[5]);
and (C[179], X[19], Y[5]);
and (C[180], X[20], Y[5]);
and (C[181], X[21], Y[5]);
and (C[182], X[22], Y[5]);
and (C[183], X[23], Y[5]);
and (C[184], X[24], Y[5]);
and (C[185], X[25], Y[5]);
and (C[186], X[26], Y[5]);
and (C[187], X[27], Y[5]);
and (C[188], X[28], Y[5]);
and (C[189], X[29], Y[5]);
and (C[190], X[30], Y[5]);
and (C[191], X[31], Y[5]);

//PP6
and (C[192], X[0], Y[6]);
and (C[193], X[1], Y[6]);
and (C[194], X[2], Y[6]);
and (C[195], X[3], Y[6]);
and (C[196], X[4], Y[6]);
and (C[197], X[5], Y[6]);
and (C[198], X[6], Y[6]);
and (C[199], X[7], Y[6]);
and (C[200], X[8], Y[6]);
and (C[201], X[9], Y[6]);
and (C[202], X[10], Y[6]);
and (C[203], X[11], Y[6]);
and (C[204], X[12], Y[6]);
and (C[205], X[13], Y[6]);
and (C[206], X[14], Y[6]);
and (C[207], X[15], Y[6]);
and (C[208], X[16], Y[6]);
and (C[209], X[17], Y[6]);
and (C[210], X[18], Y[6]);
and (C[211], X[19], Y[6]);
and (C[212], X[20], Y[6]);
and (C[213], X[21], Y[6]);
and (C[214], X[22], Y[6]);
and (C[215], X[23], Y[6]);
and (C[216], X[24], Y[6]);
and (C[217], X[25], Y[6]);
and (C[218], X[26], Y[6]);
and (C[219], X[27], Y[6]);
and (C[220], X[28], Y[6]);
and (C[221], X[29], Y[6]);
and (C[222], X[30], Y[6]);
and (C[223], X[31], Y[6]);

//PP7
and (C[224], X[0], Y[7]);
and (C[225], X[1], Y[7]);
and (C[226], X[2], Y[7]);
and (C[227], X[3], Y[7]);
and (C[228], X[4], Y[7]);
and (C[229], X[5], Y[7]);
and (C[230], X[6], Y[7]);
and (C[231], X[7], Y[7]);
and (C[232], X[8], Y[7]);
and (C[233], X[9], Y[7]);
and (C[234], X[10], Y[7]);
and (C[235], X[11], Y[7]);
and (C[236], X[12], Y[7]);
and (C[237], X[13], Y[7]);
and (C[238], X[14], Y[7]);
and (C[239], X[15], Y[7]);
and (C[240], X[16], Y[7]);
and (C[241], X[17], Y[7]);
and (C[242], X[18], Y[7]);
and (C[243], X[19], Y[7]);
and (C[244], X[20], Y[7]);
and (C[245], X[21], Y[7]);
and (C[246], X[22], Y[7]);
and (C[247], X[23], Y[7]);
and (C[248], X[24], Y[7]);
and (C[249], X[25], Y[7]);
and (C[250], X[26], Y[7]);
and (C[251], X[27], Y[7]);
and (C[252], X[28], Y[7]);
and (C[253], X[29], Y[7]);
and (C[254], X[30], Y[7]);
and (C[255], X[31], Y[7]);

//PP8
and (C[256], X[0], Y[8]);
and (C[257], X[1], Y[8]);
and (C[258], X[2], Y[8]);
and (C[259], X[3], Y[8]);
and (C[260], X[4], Y[8]);
and (C[261], X[5], Y[8]);
and (C[262], X[6], Y[8]);
and (C[263], X[7], Y[8]);
and (C[264], X[8], Y[8]);
and (C[265], X[9], Y[8]);
and (C[266], X[10], Y[8]);
and (C[267], X[11], Y[8]);
and (C[268], X[12], Y[8]);
and (C[269], X[13], Y[8]);
and (C[270], X[14], Y[8]);
and (C[271], X[15], Y[8]);
and (C[272], X[16], Y[8]);
and (C[273], X[17], Y[8]);
and (C[274], X[18], Y[8]);
and (C[275], X[19], Y[8]);
and (C[276], X[20], Y[8]);
and (C[277], X[21], Y[8]);
and (C[278], X[22], Y[8]);
and (C[279], X[23], Y[8]);
and (C[280], X[24], Y[8]);
and (C[281], X[25], Y[8]);
and (C[282], X[26], Y[8]);
and (C[283], X[27], Y[8]);
and (C[284], X[28], Y[8]);
and (C[285], X[29], Y[8]);
and (C[286], X[30], Y[8]);
and (C[287], X[31], Y[8]);

//PP9
and (C[288], X[0], Y[9]);
and (C[289], X[1], Y[9]);
and (C[290], X[2], Y[9]);
and (C[291], X[3], Y[9]);
and (C[292], X[4], Y[9]);
and (C[293], X[5], Y[9]);
and (C[294], X[6], Y[9]);
and (C[295], X[7], Y[9]);
and (C[296], X[8], Y[9]);
and (C[297], X[9], Y[9]);
and (C[298], X[10], Y[9]);
and (C[299], X[11], Y[9]);
and (C[300], X[12], Y[9]);
and (C[301], X[13], Y[9]);
and (C[302], X[14], Y[9]);
and (C[303], X[15], Y[9]);
and (C[304], X[16], Y[9]);
and (C[305], X[17], Y[9]);
and (C[306], X[18], Y[9]);
and (C[307], X[19], Y[9]);
and (C[308], X[20], Y[9]);
and (C[309], X[21], Y[9]);
and (C[310], X[22], Y[9]);
and (C[311], X[23], Y[9]);
and (C[312], X[24], Y[9]);
and (C[313], X[25], Y[9]);
and (C[314], X[26], Y[9]);
and (C[315], X[27], Y[9]);
and (C[316], X[28], Y[9]);
and (C[317], X[29], Y[9]);
and (C[318], X[30], Y[9]);
and (C[319], X[31], Y[9]);

//PP10
and (C[320], X[0], Y[10]);
and (C[321], X[1], Y[10]);
and (C[322], X[2], Y[10]);
and (C[323], X[3], Y[10]);
and (C[324], X[4], Y[10]);
and (C[325], X[5], Y[10]);
and (C[326], X[6], Y[10]);
and (C[327], X[7], Y[10]);
and (C[328], X[8], Y[10]);
and (C[329], X[9], Y[10]);
and (C[330], X[10], Y[10]);
and (C[331], X[11], Y[10]);
and (C[332], X[12], Y[10]);
and (C[333], X[13], Y[10]);
and (C[334], X[14], Y[10]);
and (C[335], X[15], Y[10]);
and (C[336], X[16], Y[10]);
and (C[337], X[17], Y[10]);
and (C[338], X[18], Y[10]);
and (C[339], X[19], Y[10]);
and (C[340], X[20], Y[10]);
and (C[341], X[21], Y[10]);
and (C[342], X[22], Y[10]);
and (C[343], X[23], Y[10]);
and (C[344], X[24], Y[10]);
and (C[345], X[25], Y[10]);
and (C[346], X[26], Y[10]);
and (C[347], X[27], Y[10]);
and (C[348], X[28], Y[10]);
and (C[349], X[29], Y[10]);
and (C[350], X[30], Y[10]);
and (C[351], X[31], Y[10]);

//PP11
and (C[352], X[0], Y[11]);
and (C[353], X[1], Y[11]);
and (C[354], X[2], Y[11]);
and (C[355], X[3], Y[11]);
and (C[356], X[4], Y[11]);
and (C[357], X[5], Y[11]);
and (C[358], X[6], Y[11]);
and (C[359], X[7], Y[11]);
and (C[360], X[8], Y[11]);
and (C[361], X[9], Y[11]);
and (C[362], X[10], Y[11]);
and (C[363], X[11], Y[11]);
and (C[364], X[12], Y[11]);
and (C[365], X[13], Y[11]);
and (C[366], X[14], Y[11]);
and (C[367], X[15], Y[11]);
and (C[368], X[16], Y[11]);
and (C[369], X[17], Y[11]);
and (C[370], X[18], Y[11]);
and (C[371], X[19], Y[11]);
and (C[372], X[20], Y[11]);
and (C[373], X[21], Y[11]);
and (C[374], X[22], Y[11]);
and (C[375], X[23], Y[11]);
and (C[376], X[24], Y[11]);
and (C[377], X[25], Y[11]);
and (C[378], X[26], Y[11]);
and (C[379], X[27], Y[11]);
and (C[380], X[28], Y[11]);
and (C[381], X[29], Y[11]);
and (C[382], X[30], Y[11]);
and (C[383], X[31], Y[11]);

//PP12
and (C[384], X[0], Y[12]);
and (C[385], X[1], Y[12]);
and (C[386], X[2], Y[12]);
and (C[387], X[3], Y[12]);
and (C[388], X[4], Y[12]);
and (C[389], X[5], Y[12]);
and (C[390], X[6], Y[12]);
and (C[391], X[7], Y[12]);
and (C[392], X[8], Y[12]);
and (C[393], X[9], Y[12]);
and (C[394], X[10], Y[12]);
and (C[395], X[11], Y[12]);
and (C[396], X[12], Y[12]);
and (C[397], X[13], Y[12]);
and (C[398], X[14], Y[12]);
and (C[399], X[15], Y[12]);
and (C[400], X[16], Y[12]);
and (C[401], X[17], Y[12]);
and (C[402], X[18], Y[12]);
and (C[403], X[19], Y[12]);
and (C[404], X[20], Y[12]);
and (C[405], X[21], Y[12]);
and (C[406], X[22], Y[12]);
and (C[407], X[23], Y[12]);
and (C[408], X[24], Y[12]);
and (C[409], X[25], Y[12]);
and (C[410], X[26], Y[12]);
and (C[411], X[27], Y[12]);
and (C[412], X[28], Y[12]);
and (C[413], X[29], Y[12]);
and (C[414], X[30], Y[12]);
and (C[415], X[31], Y[12]);

//PP13
and (C[416], X[0], Y[13]);
and (C[417], X[1], Y[13]);
and (C[418], X[2], Y[13]);
and (C[419], X[3], Y[13]);
and (C[420], X[4], Y[13]);
and (C[421], X[5], Y[13]);
and (C[422], X[6], Y[13]);
and (C[423], X[7], Y[13]);
and (C[424], X[8], Y[13]);
and (C[425], X[9], Y[13]);
and (C[426], X[10], Y[13]);
and (C[427], X[11], Y[13]);
and (C[428], X[12], Y[13]);
and (C[429], X[13], Y[13]);
and (C[430], X[14], Y[13]);
and (C[431], X[15], Y[13]);
and (C[432], X[16], Y[13]);
and (C[433], X[17], Y[13]);
and (C[434], X[18], Y[13]);
and (C[435], X[19], Y[13]);
and (C[436], X[20], Y[13]);
and (C[437], X[21], Y[13]);
and (C[438], X[22], Y[13]);
and (C[439], X[23], Y[13]);
and (C[440], X[24], Y[13]);
and (C[441], X[25], Y[13]);
and (C[442], X[26], Y[13]);
and (C[443], X[27], Y[13]);
and (C[444], X[28], Y[13]);
and (C[445], X[29], Y[13]);
and (C[446], X[30], Y[13]);
and (C[447], X[31], Y[13]);

//PP14
and (C[448], X[0], Y[14]);
and (C[449], X[1], Y[14]);
and (C[450], X[2], Y[14]);
and (C[451], X[3], Y[14]);
and (C[452], X[4], Y[14]);
and (C[453], X[5], Y[14]);
and (C[454], X[6], Y[14]);
and (C[455], X[7], Y[14]);
and (C[456], X[8], Y[14]);
and (C[457], X[9], Y[14]);
and (C[458], X[10], Y[14]);
and (C[459], X[11], Y[14]);
and (C[460], X[12], Y[14]);
and (C[461], X[13], Y[14]);
and (C[462], X[14], Y[14]);
and (C[463], X[15], Y[14]);
and (C[464], X[16], Y[14]);
and (C[465], X[17], Y[14]);
and (C[466], X[18], Y[14]);
and (C[467], X[19], Y[14]);
and (C[468], X[20], Y[14]);
and (C[469], X[21], Y[14]);
and (C[470], X[22], Y[14]);
and (C[471], X[23], Y[14]);
and (C[472], X[24], Y[14]);
and (C[473], X[25], Y[14]);
and (C[474], X[26], Y[14]);
and (C[475], X[27], Y[14]);
and (C[476], X[28], Y[14]);
and (C[477], X[29], Y[14]);
and (C[478], X[30], Y[14]);
and (C[479], X[31], Y[14]);

//PP15
and (C[480], X[0], Y[15]);
and (C[481], X[1], Y[15]);
and (C[482], X[2], Y[15]);
and (C[483], X[3], Y[15]);
and (C[484], X[4], Y[15]);
and (C[485], X[5], Y[15]);
and (C[486], X[6], Y[15]);
and (C[487], X[7], Y[15]);
and (C[488], X[8], Y[15]);
and (C[489], X[9], Y[15]);
and (C[490], X[10], Y[15]);
and (C[491], X[11], Y[15]);
and (C[492], X[12], Y[15]);
and (C[493], X[13], Y[15]);
and (C[494], X[14], Y[15]);
and (C[495], X[15], Y[15]);
and (C[496], X[16], Y[15]);
and (C[497], X[17], Y[15]);
and (C[498], X[18], Y[15]);
and (C[499], X[19], Y[15]);
and (C[500], X[20], Y[15]);
and (C[501], X[21], Y[15]);
and (C[502], X[22], Y[15]);
and (C[503], X[23], Y[15]);
and (C[504], X[24], Y[15]);
and (C[505], X[25], Y[15]);
and (C[506], X[26], Y[15]);
and (C[507], X[27], Y[15]);
and (C[508], X[28], Y[15]);
and (C[509], X[29], Y[15]);
and (C[510], X[30], Y[15]);
and (C[511], X[31], Y[15]);

//PP16
and (C[512], X[0], Y[16]);
and (C[513], X[1], Y[16]);
and (C[514], X[2], Y[16]);
and (C[515], X[3], Y[16]);
and (C[516], X[4], Y[16]);
and (C[517], X[5], Y[16]);
and (C[518], X[6], Y[16]);
and (C[519], X[7], Y[16]);
and (C[520], X[8], Y[16]);
and (C[521], X[9], Y[16]);
and (C[522], X[10], Y[16]);
and (C[523], X[11], Y[16]);
and (C[524], X[12], Y[16]);
and (C[525], X[13], Y[16]);
and (C[526], X[14], Y[16]);
and (C[527], X[15], Y[16]);
and (C[528], X[16], Y[16]);
and (C[529], X[17], Y[16]);
and (C[530], X[18], Y[16]);
and (C[531], X[19], Y[16]);
and (C[532], X[20], Y[16]);
and (C[533], X[21], Y[16]);
and (C[534], X[22], Y[16]);
and (C[535], X[23], Y[16]);
and (C[536], X[24], Y[16]);
and (C[537], X[25], Y[16]);
and (C[538], X[26], Y[16]);
and (C[539], X[27], Y[16]);
and (C[540], X[28], Y[16]);
and (C[541], X[29], Y[16]);
and (C[542], X[30], Y[16]);
and (C[543], X[31], Y[16]);

//PP17
and (C[544], X[0], Y[17]);
and (C[545], X[1], Y[17]);
and (C[546], X[2], Y[17]);
and (C[547], X[3], Y[17]);
and (C[548], X[4], Y[17]);
and (C[549], X[5], Y[17]);
and (C[550], X[6], Y[17]);
and (C[551], X[7], Y[17]);
and (C[552], X[8], Y[17]);
and (C[553], X[9], Y[17]);
and (C[554], X[10], Y[17]);
and (C[555], X[11], Y[17]);
and (C[556], X[12], Y[17]);
and (C[557], X[13], Y[17]);
and (C[558], X[14], Y[17]);
and (C[559], X[15], Y[17]);
and (C[560], X[16], Y[17]);
and (C[561], X[17], Y[17]);
and (C[562], X[18], Y[17]);
and (C[563], X[19], Y[17]);
and (C[564], X[20], Y[17]);
and (C[565], X[21], Y[17]);
and (C[566], X[22], Y[17]);
and (C[567], X[23], Y[17]);
and (C[568], X[24], Y[17]);
and (C[569], X[25], Y[17]);
and (C[570], X[26], Y[17]);
and (C[571], X[27], Y[17]);
and (C[572], X[28], Y[17]);
and (C[573], X[29], Y[17]);
and (C[574], X[30], Y[17]);
and (C[575], X[31], Y[17]);

//PP18
and (C[576], X[0], Y[18]);
and (C[577], X[1], Y[18]);
and (C[578], X[2], Y[18]);
and (C[579], X[3], Y[18]);
and (C[580], X[4], Y[18]);
and (C[581], X[5], Y[18]);
and (C[582], X[6], Y[18]);
and (C[583], X[7], Y[18]);
and (C[584], X[8], Y[18]);
and (C[585], X[9], Y[18]);
and (C[586], X[10], Y[18]);
and (C[587], X[11], Y[18]);
and (C[588], X[12], Y[18]);
and (C[589], X[13], Y[18]);
and (C[590], X[14], Y[18]);
and (C[591], X[15], Y[18]);
and (C[592], X[16], Y[18]);
and (C[593], X[17], Y[18]);
and (C[594], X[18], Y[18]);
and (C[595], X[19], Y[18]);
and (C[596], X[20], Y[18]);
and (C[597], X[21], Y[18]);
and (C[598], X[22], Y[18]);
and (C[599], X[23], Y[18]);
and (C[600], X[24], Y[18]);
and (C[601], X[25], Y[18]);
and (C[602], X[26], Y[18]);
and (C[603], X[27], Y[18]);
and (C[604], X[28], Y[18]);
and (C[605], X[29], Y[18]);
and (C[606], X[30], Y[18]);
and (C[607], X[31], Y[18]);

//PP19
and (C[608], X[0], Y[19]);
and (C[609], X[1], Y[19]);
and (C[610], X[2], Y[19]);
and (C[611], X[3], Y[19]);
and (C[612], X[4], Y[19]);
and (C[613], X[5], Y[19]);
and (C[614], X[6], Y[19]);
and (C[615], X[7], Y[19]);
and (C[616], X[8], Y[19]);
and (C[617], X[9], Y[19]);
and (C[618], X[10], Y[19]);
and (C[619], X[11], Y[19]);
and (C[620], X[12], Y[19]);
and (C[621], X[13], Y[19]);
and (C[622], X[14], Y[19]);
and (C[623], X[15], Y[19]);
and (C[624], X[16], Y[19]);
and (C[625], X[17], Y[19]);
and (C[626], X[18], Y[19]);
and (C[627], X[19], Y[19]);
and (C[628], X[20], Y[19]);
and (C[629], X[21], Y[19]);
and (C[630], X[22], Y[19]);
and (C[631], X[23], Y[19]);
and (C[632], X[24], Y[19]);
and (C[633], X[25], Y[19]);
and (C[634], X[26], Y[19]);
and (C[635], X[27], Y[19]);
and (C[636], X[28], Y[19]);
and (C[637], X[29], Y[19]);
and (C[638], X[30], Y[19]);
and (C[639], X[31], Y[19]);

//PP20
and (C[640], X[0], Y[20]);
and (C[641], X[1], Y[20]);
and (C[642], X[2], Y[20]);
and (C[643], X[3], Y[20]);
and (C[644], X[4], Y[20]);
and (C[645], X[5], Y[20]);
and (C[646], X[6], Y[20]);
and (C[647], X[7], Y[20]);
and (C[648], X[8], Y[20]);
and (C[649], X[9], Y[20]);
and (C[650], X[10], Y[20]);
and (C[651], X[11], Y[20]);
and (C[652], X[12], Y[20]);
and (C[653], X[13], Y[20]);
and (C[654], X[14], Y[20]);
and (C[655], X[15], Y[20]);
and (C[656], X[16], Y[20]);
and (C[657], X[17], Y[20]);
and (C[658], X[18], Y[20]);
and (C[659], X[19], Y[20]);
and (C[660], X[20], Y[20]);
and (C[661], X[21], Y[20]);
and (C[662], X[22], Y[20]);
and (C[663], X[23], Y[20]);
and (C[664], X[24], Y[20]);
and (C[665], X[25], Y[20]);
and (C[666], X[26], Y[20]);
and (C[667], X[27], Y[20]);
and (C[668], X[28], Y[20]);
and (C[669], X[29], Y[20]);
and (C[670], X[30], Y[20]);
and (C[671], X[31], Y[20]);

//PP21
and (C[672], X[0], Y[21]);
and (C[673], X[1], Y[21]);
and (C[674], X[2], Y[21]);
and (C[675], X[3], Y[21]);
and (C[676], X[4], Y[21]);
and (C[677], X[5], Y[21]);
and (C[678], X[6], Y[21]);
and (C[679], X[7], Y[21]);
and (C[680], X[8], Y[21]);
and (C[681], X[9], Y[21]);
and (C[682], X[10], Y[21]);
and (C[683], X[11], Y[21]);
and (C[684], X[12], Y[21]);
and (C[685], X[13], Y[21]);
and (C[686], X[14], Y[21]);
and (C[687], X[15], Y[21]);
and (C[688], X[16], Y[21]);
and (C[689], X[17], Y[21]);
and (C[690], X[18], Y[21]);
and (C[691], X[19], Y[21]);
and (C[692], X[20], Y[21]);
and (C[693], X[21], Y[21]);
and (C[694], X[22], Y[21]);
and (C[695], X[23], Y[21]);
and (C[696], X[24], Y[21]);
and (C[697], X[25], Y[21]);
and (C[698], X[26], Y[21]);
and (C[699], X[27], Y[21]);
and (C[700], X[28], Y[21]);
and (C[701], X[29], Y[21]);
and (C[702], X[30], Y[21]);
and (C[703], X[31], Y[21]);

//PP22
and (C[704], X[0], Y[22]);
and (C[705], X[1], Y[22]);
and (C[706], X[2], Y[22]);
and (C[707], X[3], Y[22]);
and (C[708], X[4], Y[22]);
and (C[709], X[5], Y[22]);
and (C[710], X[6], Y[22]);
and (C[711], X[7], Y[22]);
and (C[712], X[8], Y[22]);
and (C[713], X[9], Y[22]);
and (C[714], X[10], Y[22]);
and (C[715], X[11], Y[22]);
and (C[716], X[12], Y[22]);
and (C[717], X[13], Y[22]);
and (C[718], X[14], Y[22]);
and (C[719], X[15], Y[22]);
and (C[720], X[16], Y[22]);
and (C[721], X[17], Y[22]);
and (C[722], X[18], Y[22]);
and (C[723], X[19], Y[22]);
and (C[724], X[20], Y[22]);
and (C[725], X[21], Y[22]);
and (C[726], X[22], Y[22]);
and (C[727], X[23], Y[22]);
and (C[728], X[24], Y[22]);
and (C[729], X[25], Y[22]);
and (C[730], X[26], Y[22]);
and (C[731], X[27], Y[22]);
and (C[732], X[28], Y[22]);
and (C[733], X[29], Y[22]);
and (C[734], X[30], Y[22]);
and (C[735], X[31], Y[22]);

//PP23
and (C[736], X[0], Y[23]);
and (C[737], X[1], Y[23]);
and (C[738], X[2], Y[23]);
and (C[739], X[3], Y[23]);
and (C[740], X[4], Y[23]);
and (C[741], X[5], Y[23]);
and (C[742], X[6], Y[23]);
and (C[743], X[7], Y[23]);
and (C[744], X[8], Y[23]);
and (C[745], X[9], Y[23]);
and (C[746], X[10], Y[23]);
and (C[747], X[11], Y[23]);
and (C[748], X[12], Y[23]);
and (C[749], X[13], Y[23]);
and (C[750], X[14], Y[23]);
and (C[751], X[15], Y[23]);
and (C[752], X[16], Y[23]);
and (C[753], X[17], Y[23]);
and (C[754], X[18], Y[23]);
and (C[755], X[19], Y[23]);
and (C[756], X[20], Y[23]);
and (C[757], X[21], Y[23]);
and (C[758], X[22], Y[23]);
and (C[759], X[23], Y[23]);
and (C[760], X[24], Y[23]);
and (C[761], X[25], Y[23]);
and (C[762], X[26], Y[23]);
and (C[763], X[27], Y[23]);
and (C[764], X[28], Y[23]);
and (C[765], X[29], Y[23]);
and (C[766], X[30], Y[23]);
and (C[767], X[31], Y[23]);

//PP24
and (C[768], X[0], Y[24]);
and (C[769], X[1], Y[24]);
and (C[770], X[2], Y[24]);
and (C[771], X[3], Y[24]);
and (C[772], X[4], Y[24]);
and (C[773], X[5], Y[24]);
and (C[774], X[6], Y[24]);
and (C[775], X[7], Y[24]);
and (C[776], X[8], Y[24]);
and (C[777], X[9], Y[24]);
and (C[778], X[10], Y[24]);
and (C[779], X[11], Y[24]);
and (C[780], X[12], Y[24]);
and (C[781], X[13], Y[24]);
and (C[782], X[14], Y[24]);
and (C[783], X[15], Y[24]);
and (C[784], X[16], Y[24]);
and (C[785], X[17], Y[24]);
and (C[786], X[18], Y[24]);
and (C[787], X[19], Y[24]);
and (C[788], X[20], Y[24]);
and (C[789], X[21], Y[24]);
and (C[790], X[22], Y[24]);
and (C[791], X[23], Y[24]);
and (C[792], X[24], Y[24]);
and (C[793], X[25], Y[24]);
and (C[794], X[26], Y[24]);
and (C[795], X[27], Y[24]);
and (C[796], X[28], Y[24]);
and (C[797], X[29], Y[24]);
and (C[798], X[30], Y[24]);
and (C[799], X[31], Y[24]);

//PP25
and (C[800], X[0], Y[25]);
and (C[801], X[1], Y[25]);
and (C[802], X[2], Y[25]);
and (C[803], X[3], Y[25]);
and (C[804], X[4], Y[25]);
and (C[805], X[5], Y[25]);
and (C[806], X[6], Y[25]);
and (C[807], X[7], Y[25]);
and (C[808], X[8], Y[25]);
and (C[809], X[9], Y[25]);
and (C[810], X[10], Y[25]);
and (C[811], X[11], Y[25]);
and (C[812], X[12], Y[25]);
and (C[813], X[13], Y[25]);
and (C[814], X[14], Y[25]);
and (C[815], X[15], Y[25]);
and (C[816], X[16], Y[25]);
and (C[817], X[17], Y[25]);
and (C[818], X[18], Y[25]);
and (C[819], X[19], Y[25]);
and (C[820], X[20], Y[25]);
and (C[821], X[21], Y[25]);
and (C[822], X[22], Y[25]);
and (C[823], X[23], Y[25]);
and (C[824], X[24], Y[25]);
and (C[825], X[25], Y[25]);
and (C[826], X[26], Y[25]);
and (C[827], X[27], Y[25]);
and (C[828], X[28], Y[25]);
and (C[829], X[29], Y[25]);
and (C[830], X[30], Y[25]);
and (C[831], X[31], Y[25]);

//PP26
and (C[832], X[0], Y[26]);
and (C[833], X[1], Y[26]);
and (C[834], X[2], Y[26]);
and (C[835], X[3], Y[26]);
and (C[836], X[4], Y[26]);
and (C[837], X[5], Y[26]);
and (C[838], X[6], Y[26]);
and (C[839], X[7], Y[26]);
and (C[840], X[8], Y[26]);
and (C[841], X[9], Y[26]);
and (C[842], X[10], Y[26]);
and (C[843], X[11], Y[26]);
and (C[844], X[12], Y[26]);
and (C[845], X[13], Y[26]);
and (C[846], X[14], Y[26]);
and (C[847], X[15], Y[26]);
and (C[848], X[16], Y[26]);
and (C[849], X[17], Y[26]);
and (C[850], X[18], Y[26]);
and (C[851], X[19], Y[26]);
and (C[852], X[20], Y[26]);
and (C[853], X[21], Y[26]);
and (C[854], X[22], Y[26]);
and (C[855], X[23], Y[26]);
and (C[856], X[24], Y[26]);
and (C[857], X[25], Y[26]);
and (C[858], X[26], Y[26]);
and (C[859], X[27], Y[26]);
and (C[860], X[28], Y[26]);
and (C[861], X[29], Y[26]);
and (C[862], X[30], Y[26]);
and (C[863], X[31], Y[26]);

//PP27
and (C[864], X[0], Y[27]);
and (C[865], X[1], Y[27]);
and (C[866], X[2], Y[27]);
and (C[867], X[3], Y[27]);
and (C[868], X[4], Y[27]);
and (C[869], X[5], Y[27]);
and (C[870], X[6], Y[27]);
and (C[871], X[7], Y[27]);
and (C[872], X[8], Y[27]);
and (C[873], X[9], Y[27]);
and (C[874], X[10], Y[27]);
and (C[875], X[11], Y[27]);
and (C[876], X[12], Y[27]);
and (C[877], X[13], Y[27]);
and (C[878], X[14], Y[27]);
and (C[879], X[15], Y[27]);
and (C[880], X[16], Y[27]);
and (C[881], X[17], Y[27]);
and (C[882], X[18], Y[27]);
and (C[883], X[19], Y[27]);
and (C[884], X[20], Y[27]);
and (C[885], X[21], Y[27]);
and (C[886], X[22], Y[27]);
and (C[887], X[23], Y[27]);
and (C[888], X[24], Y[27]);
and (C[889], X[25], Y[27]);
and (C[890], X[26], Y[27]);
and (C[891], X[27], Y[27]);
and (C[892], X[28], Y[27]);
and (C[893], X[29], Y[27]);
and (C[894], X[30], Y[27]);
and (C[895], X[31], Y[27]);

//PP28
and (C[896], X[0], Y[28]);
and (C[897], X[1], Y[28]);
and (C[898], X[2], Y[28]);
and (C[899], X[3], Y[28]);
and (C[900], X[4], Y[28]);
and (C[901], X[5], Y[28]);
and (C[902], X[6], Y[28]);
and (C[903], X[7], Y[28]);
and (C[904], X[8], Y[28]);
and (C[905], X[9], Y[28]);
and (C[906], X[10], Y[28]);
and (C[907], X[11], Y[28]);
and (C[908], X[12], Y[28]);
and (C[909], X[13], Y[28]);
and (C[910], X[14], Y[28]);
and (C[911], X[15], Y[28]);
and (C[912], X[16], Y[28]);
and (C[913], X[17], Y[28]);
and (C[914], X[18], Y[28]);
and (C[915], X[19], Y[28]);
and (C[916], X[20], Y[28]);
and (C[917], X[21], Y[28]);
and (C[918], X[22], Y[28]);
and (C[919], X[23], Y[28]);
and (C[920], X[24], Y[28]);
and (C[921], X[25], Y[28]);
and (C[922], X[26], Y[28]);
and (C[923], X[27], Y[28]);
and (C[924], X[28], Y[28]);
and (C[925], X[29], Y[28]);
and (C[926], X[30], Y[28]);
and (C[927], X[31], Y[28]);

//PP29
and (C[928], X[0], Y[29]);
and (C[929], X[1], Y[29]);
and (C[930], X[2], Y[29]);
and (C[931], X[3], Y[29]);
and (C[932], X[4], Y[29]);
and (C[933], X[5], Y[29]);
and (C[934], X[6], Y[29]);
and (C[935], X[7], Y[29]);
and (C[936], X[8], Y[29]);
and (C[937], X[9], Y[29]);
and (C[938], X[10], Y[29]);
and (C[939], X[11], Y[29]);
and (C[940], X[12], Y[29]);
and (C[941], X[13], Y[29]);
and (C[942], X[14], Y[29]);
and (C[943], X[15], Y[29]);
and (C[944], X[16], Y[29]);
and (C[945], X[17], Y[29]);
and (C[946], X[18], Y[29]);
and (C[947], X[19], Y[29]);
and (C[948], X[20], Y[29]);
and (C[949], X[21], Y[29]);
and (C[950], X[22], Y[29]);
and (C[951], X[23], Y[29]);
and (C[952], X[24], Y[29]);
and (C[953], X[25], Y[29]);
and (C[954], X[26], Y[29]);
and (C[955], X[27], Y[29]);
and (C[956], X[28], Y[29]);
and (C[957], X[29], Y[29]);
and (C[958], X[30], Y[29]);
and (C[959], X[31], Y[29]);

//PP30
and (C[960], X[0], Y[30]);
and (C[961], X[1], Y[30]);
and (C[962], X[2], Y[30]);
and (C[963], X[3], Y[30]);
and (C[964], X[4], Y[30]);
and (C[965], X[5], Y[30]);
and (C[966], X[6], Y[30]);
and (C[967], X[7], Y[30]);
and (C[968], X[8], Y[30]);
and (C[969], X[9], Y[30]);
and (C[970], X[10], Y[30]);
and (C[971], X[11], Y[30]);
and (C[972], X[12], Y[30]);
and (C[973], X[13], Y[30]);
and (C[974], X[14], Y[30]);
and (C[975], X[15], Y[30]);
and (C[976], X[16], Y[30]);
and (C[977], X[17], Y[30]);
and (C[978], X[18], Y[30]);
and (C[979], X[19], Y[30]);
and (C[980], X[20], Y[30]);
and (C[981], X[21], Y[30]);
and (C[982], X[22], Y[30]);
and (C[983], X[23], Y[30]);
and (C[984], X[24], Y[30]);
and (C[985], X[25], Y[30]);
and (C[986], X[26], Y[30]);
and (C[987], X[27], Y[30]);
and (C[988], X[28], Y[30]);
and (C[989], X[29], Y[30]);
and (C[990], X[30], Y[30]);
and (C[991], X[31], Y[30]);

//PP31
and (C[992], X[0], Y[31]);
and (C[993], X[1], Y[31]);
and (C[994], X[2], Y[31]);
and (C[995], X[3], Y[31]);
and (C[996], X[4], Y[31]);
and (C[997], X[5], Y[31]);
and (C[998], X[6], Y[31]);
and (C[999], X[7], Y[31]);
and (C[1000], X[8], Y[31]);
and (C[1001], X[9], Y[31]);
and (C[1002], X[10], Y[31]);
and (C[1003], X[11], Y[31]);
and (C[1004], X[12], Y[31]);
and (C[1005], X[13], Y[31]);
and (C[1006], X[14], Y[31]);
and (C[1007], X[15], Y[31]);
and (C[1008], X[16], Y[31]);
and (C[1009], X[17], Y[31]);
and (C[1010], X[18], Y[31]);
and (C[1011], X[19], Y[31]);
and (C[1012], X[20], Y[31]);
and (C[1013], X[21], Y[31]);
and (C[1014], X[22], Y[31]);
and (C[1015], X[23], Y[31]);
and (C[1016], X[24], Y[31]);
and (C[1017], X[25], Y[31]);
and (C[1018], X[26], Y[31]);
and (C[1019], X[27], Y[31]);
and (C[1020], X[28], Y[31]);
and (C[1021], X[29], Y[31]);
and (C[1022], X[30], Y[31]);
and (C[1023], X[31], Y[31]);


//pp0,1,2
fulladd full00(sum[0], carry[0], C[0], 1'b0, 1'b0);
fulladd full01(sum[1], carry[1], C[1], C[32], 1'b0);
fulladd full02 (sum[2], carry[2], C[2], C[33], C[64] );
fulladd full03 (sum[3], carry[3], C[3], C[34], C[65] );
fulladd full04 (sum[4], carry[4], C[4], C[35], C[66] );
fulladd full05 (sum[5], carry[5], C[5], C[36], C[67] );
fulladd full06 (sum[6], carry[6], C[6], C[37], C[68] );
fulladd full07 (sum[7], carry[7], C[7], C[38], C[69] );
fulladd full08 (sum[8], carry[8], C[8], C[39], C[70] );
fulladd full09 (sum[9], carry[9], C[9], C[40], C[71] );
fulladd full010 (sum[10], carry[10], C[10], C[41], C[72] );
fulladd full011 (sum[11], carry[11], C[11], C[42], C[73] );
fulladd full012 (sum[12], carry[12], C[12], C[43], C[74] );
fulladd full013 (sum[13], carry[13], C[13], C[44], C[75] );
fulladd full014 (sum[14], carry[14], C[14], C[45], C[76] );
fulladd full015 (sum[15], carry[15], C[15], C[46], C[77] );
fulladd full016 (sum[16], carry[16], C[16], C[47], C[78] );
fulladd full017 (sum[17], carry[17], C[17], C[48], C[79] );
fulladd full018 (sum[18], carry[18], C[18], C[49], C[80] );
fulladd full019 (sum[19], carry[19], C[19], C[50], C[81] );
fulladd full020 (sum[20], carry[20], C[20], C[51], C[82] );
fulladd full021 (sum[21], carry[21], C[21], C[52], C[83] );
fulladd full022 (sum[22], carry[22], C[22], C[53], C[84] );
fulladd full023 (sum[23], carry[23], C[23], C[54], C[85] );
fulladd full024 (sum[24], carry[24], C[24], C[55], C[86] );
fulladd full025 (sum[25], carry[25], C[25], C[56], C[87] );
fulladd full026 (sum[26], carry[26], C[26], C[57], C[88] );
fulladd full027 (sum[27], carry[27], C[27], C[58], C[89] );
fulladd full028 (sum[28], carry[28], C[28], C[59], C[90] );
fulladd full029 (sum[29], carry[29], C[29], C[60], C[91] );
fulladd full030 (sum[30], carry[30], C[30], C[61], C[92] );
fulladd full031 (sum[31], carry[31], C[31], C[62], C[93] );
fulladd full032 (sum[32], carry[32], 1'b0, C[63], C[94] );
fulladd full033 (sum[33], carry[33], 1'b0, 1'b0, C[95] );
fulladd full034 (sum[34], carry[34], 1'b0, 1'b0, 1'b0 );
fulladd full035 (sum[35], carry[35], 1'b0, 1'b0, 1'b0 );
fulladd full036 (sum[36], carry[36], 1'b0, 1'b0, 1'b0 );
fulladd full037 (sum[37], carry[37], 1'b0, 1'b0, 1'b0 );
fulladd full038 (sum[38], carry[38], 1'b0, 1'b0, 1'b0 );
fulladd full039 (sum[39], carry[39], 1'b0, 1'b0, 1'b0 );
fulladd full040 (sum[40], carry[40], 1'b0, 1'b0, 1'b0 );
fulladd full041 (sum[41], carry[41], 1'b0, 1'b0, 1'b0 );
fulladd full042 (sum[42], carry[42], 1'b0, 1'b0, 1'b0 );
fulladd full043 (sum[43], carry[43], 1'b0, 1'b0, 1'b0 );
fulladd full044 (sum[44], carry[44], 1'b0, 1'b0, 1'b0 );
fulladd full045 (sum[45], carry[45], 1'b0, 1'b0, 1'b0 );
fulladd full046 (sum[46], carry[46], 1'b0, 1'b0, 1'b0 );
fulladd full047 (sum[47], carry[47], 1'b0, 1'b0, 1'b0 );
fulladd full048 (sum[48], carry[48], 1'b0, 1'b0, 1'b0 );
fulladd full049 (sum[49], carry[49], 1'b0, 1'b0, 1'b0 );
fulladd full050 (sum[50], carry[50], 1'b0, 1'b0, 1'b0 );
fulladd full051 (sum[51], carry[51], 1'b0, 1'b0, 1'b0 );
fulladd full052 (sum[52], carry[52], 1'b0, 1'b0, 1'b0 );
fulladd full053 (sum[53], carry[53], 1'b0, 1'b0, 1'b0 );
fulladd full054 (sum[54], carry[54], 1'b0, 1'b0, 1'b0 );
fulladd full055 (sum[55], carry[55], 1'b0, 1'b0, 1'b0 );
fulladd full056 (sum[56], carry[56], 1'b0, 1'b0, 1'b0 );
fulladd full057 (sum[57], carry[57], 1'b0, 1'b0, 1'b0 );
fulladd full058 (sum[58], carry[58], 1'b0, 1'b0, 1'b0 );
fulladd full059 (sum[59], carry[59], 1'b0, 1'b0, 1'b0 );
fulladd full060 (sum[60], carry[60], 1'b0, 1'b0, 1'b0 );
fulladd full061 (sum[61], carry[61], 1'b0, 1'b0, 1'b0 );
fulladd full062 (sum[62], carry[62], 1'b0, 1'b0, 1'b0 );
fulladd full063 (sum[63], carry[63], 1'b0, 1'b0, 1'b0 );

//pp3,4,5
fulladd full10(sum[64], carry[64], 1'b0, 1'b0, 1'b0);
fulladd full11(sum[65], carry[65], 1'b0, 1'b0, 1'b0);
fulladd full12(sum[66], carry[66], 1'b0, 1'b0, 1'b0);
fulladd full13(sum[67], carry[67], C[96], 1'b0, 1'b0);
fulladd full14(sum[68], carry[68], C[97], C[128], 1'b0);
fulladd full15 (sum[69], carry[69], C[98], C[129], C[160]);
fulladd full16 (sum[70], carry[70], C[99], C[130], C[161]);
fulladd full17 (sum[71], carry[71], C[100], C[131], C[162]);
fulladd full18 (sum[72], carry[72], C[101], C[132], C[163]);
fulladd full19 (sum[73], carry[73], C[102], C[133], C[164]);
fulladd full110 (sum[74], carry[74], C[103], C[134], C[165]);
fulladd full111 (sum[75], carry[75], C[104], C[135], C[166]);
fulladd full112 (sum[76], carry[76], C[105], C[136], C[167]);
fulladd full113 (sum[77], carry[77], C[106], C[137], C[168]);
fulladd full114 (sum[78], carry[78], C[107], C[138], C[169]);
fulladd full115 (sum[79], carry[79], C[108], C[139], C[170]);
fulladd full116 (sum[80], carry[80], C[109], C[140], C[171]);
fulladd full117 (sum[81], carry[81], C[110], C[141], C[172]);
fulladd full118 (sum[82], carry[82], C[111], C[142], C[173]);
fulladd full119 (sum[83], carry[83], C[112], C[143], C[174]);
fulladd full120 (sum[84], carry[84], C[113], C[144], C[175]);
fulladd full121 (sum[85], carry[85], C[114], C[145], C[176]);
fulladd full122 (sum[86], carry[86], C[115], C[146], C[177]);
fulladd full123 (sum[87], carry[87], C[116], C[147], C[178]);
fulladd full124 (sum[88], carry[88], C[117], C[148], C[179]);
fulladd full125 (sum[89], carry[89], C[118], C[149], C[180]);
fulladd full126 (sum[90], carry[90], C[119], C[150], C[181]);
fulladd full127 (sum[91], carry[91], C[120], C[151], C[182]);
fulladd full128 (sum[92], carry[92], C[121], C[152], C[183]);
fulladd full129 (sum[93], carry[93], C[122], C[153], C[184]);
fulladd full130 (sum[94], carry[94], C[123], C[154], C[185]);
fulladd full131 (sum[95], carry[95], C[124], C[155], C[186]);
fulladd full132 (sum[96], carry[96], C[125], C[156], C[187]);
fulladd full133 (sum[97], carry[97], C[126], C[157], C[188]);
fulladd full134 (sum[98], carry[98], C[127], C[158], C[189]);
fulladd full135 (sum[99], carry[99], 1'b0, C[159], C[190]);
fulladd full136 (sum[100], carry[100], 1'b0, 1'b0, C[191]);
fulladd full137 (sum[101], carry[101], 1'b0, 1'b0, 1'b0);
fulladd full138 (sum[102], carry[102], 1'b0, 1'b0, 1'b0);
fulladd full139 (sum[103], carry[103], 1'b0, 1'b0, 1'b0);
fulladd full140 (sum[104], carry[104], 1'b0, 1'b0, 1'b0);
fulladd full141 (sum[105], carry[105], 1'b0, 1'b0, 1'b0);
fulladd full142 (sum[106], carry[106], 1'b0, 1'b0, 1'b0);
fulladd full143 (sum[107], carry[107], 1'b0, 1'b0, 1'b0);
fulladd full144 (sum[108], carry[108], 1'b0, 1'b0, 1'b0);
fulladd full145 (sum[109], carry[109], 1'b0, 1'b0, 1'b0);
fulladd full146 (sum[110], carry[110], 1'b0, 1'b0, 1'b0);
fulladd full147 (sum[111], carry[111], 1'b0, 1'b0, 1'b0);
fulladd full148 (sum[112], carry[112], 1'b0, 1'b0, 1'b0);
fulladd full149 (sum[113], carry[113], 1'b0, 1'b0, 1'b0);
fulladd full150 (sum[114], carry[114], 1'b0, 1'b0, 1'b0);
fulladd full151 (sum[115], carry[115], 1'b0, 1'b0, 1'b0);
fulladd full152 (sum[116], carry[116], 1'b0, 1'b0, 1'b0);
fulladd full153 (sum[117], carry[117], 1'b0, 1'b0, 1'b0);
fulladd full154 (sum[118], carry[118], 1'b0, 1'b0, 1'b0);
fulladd full155 (sum[119], carry[119], 1'b0, 1'b0, 1'b0);
fulladd full156 (sum[120], carry[120], 1'b0, 1'b0, 1'b0);
fulladd full157 (sum[121], carry[121], 1'b0, 1'b0, 1'b0);
fulladd full158 (sum[122], carry[122], 1'b0, 1'b0, 1'b0);
fulladd full159 (sum[123], carry[123], 1'b0, 1'b0, 1'b0);
fulladd full160 (sum[124], carry[124], 1'b0, 1'b0, 1'b0);
fulladd full161 (sum[125], carry[125], 1'b0, 1'b0, 1'b0);
fulladd full162 (sum[126], carry[126], 1'b0, 1'b0, 1'b0);
fulladd full163 (sum[127], carry[127], 1'b0, 1'b0, 1'b0);

//pp6,7,8
fulladd full20 (sum[128], carry[128], 1'b0, 1'b0, 1'b0);
fulladd full21 (sum[129], carry[129], 1'b0, 1'b0, 1'b0);
fulladd full22 (sum[130], carry[130], 1'b0, 1'b0, 1'b0);
fulladd full23 (sum[131], carry[131], 1'b0, 1'b0, 1'b0);
fulladd full24 (sum[132], carry[132], 1'b0, 1'b0, 1'b0);
fulladd full25 (sum[133], carry[133], 1'b0, 1'b0, 1'b0);
fulladd full26 (sum[134], carry[134], C[192], 1'b0, 1'b0);
fulladd full27 (sum[135], carry[135], C[193], C[224], 1'b0);
fulladd full28 (sum[136], carry[136], C[194], C[225], C[256]);
fulladd full29 (sum[137], carry[137], C[195], C[226], C[257]);
fulladd full210 (sum[138], carry[138], C[196], C[227], C[258]);
fulladd full211 (sum[139], carry[139], C[197], C[228], C[259]);
fulladd full212 (sum[140], carry[140], C[198], C[229], C[260]);
fulladd full213 (sum[141], carry[141], C[199], C[230], C[261]);
fulladd full214 (sum[142], carry[142], C[200], C[231], C[262]);
fulladd full215 (sum[143], carry[143], C[201], C[232], C[263]);
fulladd full216 (sum[144], carry[144], C[202], C[233], C[264]);
fulladd full217 (sum[145], carry[145], C[203], C[234], C[265]);
fulladd full218 (sum[146], carry[146], C[204], C[235], C[266]);
fulladd full219 (sum[147], carry[147], C[205], C[236], C[267]);
fulladd full220 (sum[148], carry[148], C[206], C[237], C[268]);
fulladd full221 (sum[149], carry[149], C[207], C[238], C[269]);
fulladd full222 (sum[150], carry[150], C[208], C[239], C[270]);
fulladd full223 (sum[151], carry[151], C[209], C[240], C[271]);
fulladd full224 (sum[152], carry[152], C[210], C[241], C[272]);
fulladd full225 (sum[153], carry[153], C[211], C[242], C[273]);
fulladd full226 (sum[154], carry[154], C[212], C[243], C[274]);
fulladd full227 (sum[155], carry[155], C[213], C[244], C[275]);
fulladd full228 (sum[156], carry[156], C[214], C[245], C[276]);
fulladd full229 (sum[157], carry[157], C[215], C[246], C[277]);
fulladd full230 (sum[158], carry[158], C[216], C[247], C[278]);
fulladd full231 (sum[159], carry[159], C[217], C[248], C[279]);
fulladd full232 (sum[160], carry[160], C[218], C[249], C[280]);
fulladd full233 (sum[161], carry[161], C[219], C[250], C[281]);
fulladd full234 (sum[162], carry[162], C[220], C[251], C[282]);
fulladd full235 (sum[163], carry[163], C[221], C[252], C[283]);
fulladd full236 (sum[164], carry[164], C[222], C[253], C[284]);
fulladd full237 (sum[165], carry[165], C[223], C[254], C[285]);
fulladd full238 (sum[166], carry[166], 1'b0, C[255], C[286]);
fulladd full239 (sum[167], carry[167], 1'b0, 1'b0, C[287]);
fulladd full240 (sum[168], carry[168], 1'b0, 1'b0, 1'b0);
fulladd full241 (sum[169], carry[169], 1'b0, 1'b0, 1'b0);
fulladd full242 (sum[170], carry[170], 1'b0, 1'b0, 1'b0);
fulladd full243 (sum[171], carry[171], 1'b0, 1'b0, 1'b0);
fulladd full244 (sum[172], carry[172], 1'b0, 1'b0, 1'b0);
fulladd full245 (sum[173], carry[173], 1'b0, 1'b0, 1'b0);
fulladd full246 (sum[174], carry[174], 1'b0, 1'b0, 1'b0);
fulladd full247 (sum[175], carry[175], 1'b0, 1'b0, 1'b0);
fulladd full248 (sum[176], carry[176], 1'b0, 1'b0, 1'b0);
fulladd full249 (sum[177], carry[177], 1'b0, 1'b0, 1'b0);
fulladd full250 (sum[178], carry[178], 1'b0, 1'b0, 1'b0);
fulladd full251 (sum[179], carry[179], 1'b0, 1'b0, 1'b0);
fulladd full252 (sum[180], carry[180], 1'b0, 1'b0, 1'b0);
fulladd full253 (sum[181], carry[181], 1'b0, 1'b0, 1'b0);
fulladd full254 (sum[182], carry[182], 1'b0, 1'b0, 1'b0);
fulladd full255 (sum[183], carry[183], 1'b0, 1'b0, 1'b0);
fulladd full256 (sum[184], carry[184], 1'b0, 1'b0, 1'b0);
fulladd full257 (sum[185], carry[185], 1'b0, 1'b0, 1'b0);
fulladd full258 (sum[186], carry[186], 1'b0, 1'b0, 1'b0);
fulladd full259 (sum[187], carry[187], 1'b0, 1'b0, 1'b0);
fulladd full260 (sum[188], carry[188], 1'b0, 1'b0, 1'b0);
fulladd full261 (sum[189], carry[189], 1'b0, 1'b0, 1'b0);
fulladd full262 (sum[190], carry[190], 1'b0, 1'b0, 1'b0);
fulladd full263 (sum[191], carry[191], 1'b0, 1'b0, 1'b0);

//pp9,10,11
fulladd full30 (sum[192], carry[192], 1'b0, 1'b0, 1'b0);
fulladd full31 (sum[193], carry[193], 1'b0, 1'b0, 1'b0);
fulladd full32 (sum[194], carry[194], 1'b0, 1'b0, 1'b0);
fulladd full33 (sum[195], carry[195], 1'b0, 1'b0, 1'b0);
fulladd full34 (sum[196], carry[196], 1'b0, 1'b0, 1'b0);
fulladd full35 (sum[197], carry[197], 1'b0, 1'b0, 1'b0);
fulladd full36 (sum[198], carry[198], 1'b0, 1'b0, 1'b0);
fulladd full37 (sum[199], carry[199], 1'b0, 1'b0, 1'b0);
fulladd full38 (sum[200], carry[200], 1'b0, 1'b0, 1'b0);
fulladd full39 (sum[201], carry[201], C[288], 1'b0, 1'b0);
fulladd full310 (sum[202], carry[202], C[289], C[320], 1'b0);
fulladd full311 (sum[203], carry[203], C[290], C[321], C[352]);
fulladd full312 (sum[204], carry[204], C[291], C[322], C[353]);
fulladd full313 (sum[205], carry[205], C[292], C[323], C[354]);
fulladd full314 (sum[206], carry[206], C[293], C[324], C[355]);
fulladd full315 (sum[207], carry[207], C[294], C[325], C[356]);
fulladd full316 (sum[208], carry[208], C[295], C[326], C[357]);
fulladd full317 (sum[209], carry[209], C[296], C[327], C[358]);
fulladd full318 (sum[210], carry[210], C[297], C[328], C[359]);
fulladd full319 (sum[211], carry[211], C[298], C[329], C[360]);
fulladd full320 (sum[212], carry[212], C[299], C[330], C[361]);
fulladd full321 (sum[213], carry[213], C[300], C[331], C[362]);
fulladd full322 (sum[214], carry[214], C[301], C[332], C[363]);
fulladd full323 (sum[215], carry[215], C[302], C[333], C[364]);
fulladd full324 (sum[216], carry[216], C[303], C[334], C[365]);
fulladd full325 (sum[217], carry[217], C[304], C[335], C[366]);
fulladd full326 (sum[218], carry[218], C[305], C[336], C[367]);
fulladd full327 (sum[219], carry[219], C[306], C[337], C[368]);
fulladd full328 (sum[220], carry[220], C[307], C[338], C[369]);
fulladd full329 (sum[221], carry[221], C[308], C[339], C[370]);
fulladd full330 (sum[222], carry[222], C[309], C[340], C[371]);
fulladd full331 (sum[223], carry[223], C[310], C[341], C[372]);
fulladd full332 (sum[224], carry[224], C[311], C[342], C[373]);
fulladd full333 (sum[225], carry[225], C[312], C[343], C[374]);
fulladd full334 (sum[226], carry[226], C[313], C[344], C[375]);
fulladd full335 (sum[227], carry[227], C[314], C[345], C[376]);
fulladd full336 (sum[228], carry[228], C[315], C[346], C[377]);
fulladd full337 (sum[229], carry[229], C[316], C[347], C[378]);
fulladd full338 (sum[230], carry[230], C[317], C[348], C[379]);
fulladd full339 (sum[231], carry[231], C[318], C[349], C[380]);
fulladd full340 (sum[232], carry[232], C[319], C[350], C[381]);
fulladd full341 (sum[233], carry[233], 1'b0, C[351], C[382]);
fulladd full342 (sum[234], carry[234], 1'b0, 1'b0, C[383]);
fulladd full343 (sum[235], carry[235], 1'b0, 1'b0, 1'b0);
fulladd full344 (sum[236], carry[236], 1'b0, 1'b0, 1'b0);
fulladd full345 (sum[237], carry[237], 1'b0, 1'b0, 1'b0);
fulladd full346 (sum[238], carry[238], 1'b0, 1'b0, 1'b0);
fulladd full347 (sum[239], carry[239], 1'b0, 1'b0, 1'b0);
fulladd full348 (sum[240], carry[240], 1'b0, 1'b0, 1'b0);
fulladd full349 (sum[241], carry[241], 1'b0, 1'b0, 1'b0);
fulladd full350 (sum[242], carry[242], 1'b0, 1'b0, 1'b0);
fulladd full351 (sum[243], carry[243], 1'b0, 1'b0, 1'b0);
fulladd full352 (sum[244], carry[244], 1'b0, 1'b0, 1'b0);
fulladd full353 (sum[245], carry[245], 1'b0, 1'b0, 1'b0);
fulladd full354 (sum[246], carry[246], 1'b0, 1'b0, 1'b0);
fulladd full355 (sum[247], carry[247], 1'b0, 1'b0, 1'b0);
fulladd full356 (sum[248], carry[248], 1'b0, 1'b0, 1'b0);
fulladd full357 (sum[249], carry[249], 1'b0, 1'b0, 1'b0);
fulladd full358 (sum[250], carry[250], 1'b0, 1'b0, 1'b0);
fulladd full359 (sum[251], carry[251], 1'b0, 1'b0, 1'b0);
fulladd full360 (sum[252], carry[252], 1'b0, 1'b0, 1'b0);
fulladd full361 (sum[253], carry[253], 1'b0, 1'b0, 1'b0);
fulladd full362 (sum[254], carry[254], 1'b0, 1'b0, 1'b0);
fulladd full363 (sum[255], carry[255], 1'b0, 1'b0, 1'b0);

//pp12,13,14
fulladd full40 (sum[256], carry[256], 1'b0, 1'b0, 1'b0);
fulladd full41 (sum[257], carry[257], 1'b0, 1'b0, 1'b0);
fulladd full42 (sum[258], carry[258], 1'b0, 1'b0, 1'b0);
fulladd full43 (sum[259], carry[259], 1'b0, 1'b0, 1'b0);
fulladd full44 (sum[260], carry[260], 1'b0, 1'b0, 1'b0);
fulladd full45 (sum[261], carry[261], 1'b0, 1'b0, 1'b0);
fulladd full46 (sum[262], carry[262], 1'b0, 1'b0, 1'b0);
fulladd full47 (sum[263], carry[263], 1'b0, 1'b0, 1'b0);
fulladd full48 (sum[264], carry[264], 1'b0, 1'b0, 1'b0);
fulladd full49 (sum[265], carry[265], 1'b0, 1'b0, 1'b0);
fulladd full410 (sum[266], carry[266], 1'b0, 1'b0, 1'b0);
fulladd full411 (sum[267], carry[267], 1'b0, 1'b0, 1'b0);
fulladd full412 (sum[268], carry[268], C[384], 1'b0, 1'b0);
fulladd full413 (sum[269], carry[269], C[385], C[416], 1'b0);
fulladd full414 (sum[270], carry[270], C[386], C[417], C[448]);
fulladd full415 (sum[271], carry[271], C[387], C[418], C[449]);
fulladd full416 (sum[272], carry[272], C[388], C[419], C[450]);
fulladd full417 (sum[273], carry[273], C[389], C[420], C[451]);
fulladd full418 (sum[274], carry[274], C[390], C[421], C[452]);
fulladd full419 (sum[275], carry[275], C[391], C[422], C[453]);
fulladd full420 (sum[276], carry[276], C[392], C[423], C[454]);
fulladd full421 (sum[277], carry[277], C[393], C[424], C[455]);
fulladd full422 (sum[278], carry[278], C[394], C[425], C[456]);
fulladd full423 (sum[279], carry[279], C[395], C[426], C[457]);
fulladd full424 (sum[280], carry[280], C[396], C[427], C[458]);
fulladd full425 (sum[281], carry[281], C[397], C[428], C[459]);
fulladd full426 (sum[282], carry[282], C[398], C[429], C[460]);
fulladd full427 (sum[283], carry[283], C[399], C[430], C[461]);
fulladd full428 (sum[284], carry[284], C[400], C[431], C[462]);
fulladd full429 (sum[285], carry[285], C[401], C[432], C[463]);
fulladd full430 (sum[286], carry[286], C[402], C[433], C[464]);
fulladd full431 (sum[287], carry[287], C[403], C[434], C[465]);
fulladd full432 (sum[288], carry[288], C[404], C[435], C[466]);
fulladd full433 (sum[289], carry[289], C[405], C[436], C[467]);
fulladd full434 (sum[290], carry[290], C[406], C[437], C[468]);
fulladd full435 (sum[291], carry[291], C[407], C[438], C[469]);
fulladd full436 (sum[292], carry[292], C[408], C[439], C[470]);
fulladd full437 (sum[293], carry[293], C[409], C[440], C[471]);
fulladd full438 (sum[294], carry[294], C[410], C[441], C[472]);
fulladd full439 (sum[295], carry[295], C[411], C[442], C[473]);
fulladd full440 (sum[296], carry[296], C[412], C[443], C[474]);
fulladd full441 (sum[297], carry[297], C[413], C[444], C[475]);
fulladd full442 (sum[298], carry[298], C[414], C[445], C[476]);
fulladd full443 (sum[299], carry[299], C[415], C[446], C[477]);
fulladd full444 (sum[300], carry[300], 1'b0, C[477], C[478]);
fulladd full445 (sum[301], carry[301], 1'b0, 1'b0, C[479]);
fulladd full446 (sum[302], carry[302], 1'b0, 1'b0, 1'b0);
fulladd full447 (sum[303], carry[303], 1'b0, 1'b0, 1'b0);
fulladd full448 (sum[304], carry[304], 1'b0, 1'b0, 1'b0);
fulladd full449 (sum[305], carry[305], 1'b0, 1'b0, 1'b0);
fulladd full450 (sum[306], carry[306], 1'b0, 1'b0, 1'b0);
fulladd full451 (sum[307], carry[307], 1'b0, 1'b0, 1'b0);
fulladd full452 (sum[308], carry[308], 1'b0, 1'b0, 1'b0);
fulladd full453 (sum[309], carry[309], 1'b0, 1'b0, 1'b0);
fulladd full454 (sum[310], carry[310], 1'b0, 1'b0, 1'b0);
fulladd full455 (sum[311], carry[311], 1'b0, 1'b0, 1'b0);
fulladd full456 (sum[312], carry[312], 1'b0, 1'b0, 1'b0);
fulladd full457 (sum[313], carry[313], 1'b0, 1'b0, 1'b0);
fulladd full458 (sum[314], carry[314], 1'b0, 1'b0, 1'b0);
fulladd full459 (sum[315], carry[315], 1'b0, 1'b0, 1'b0);
fulladd full460 (sum[316], carry[316], 1'b0, 1'b0, 1'b0);
fulladd full461 (sum[317], carry[317], 1'b0, 1'b0, 1'b0);
fulladd full462 (sum[318], carry[318], 1'b0, 1'b0, 1'b0);
fulladd full463 (sum[319], carry[319], 1'b0, 1'b0, 1'b0);

//pp15,16,17
fulladd full50 (sum[320], carry[320], 1'b0, 1'b0, 1'b0);
fulladd full51 (sum[321], carry[321], 1'b0, 1'b0, 1'b0);
fulladd full52 (sum[322], carry[322], 1'b0, 1'b0, 1'b0);
fulladd full53 (sum[323], carry[323], 1'b0, 1'b0, 1'b0);
fulladd full54 (sum[324], carry[324], 1'b0, 1'b0, 1'b0);
fulladd full55 (sum[325], carry[325], 1'b0, 1'b0, 1'b0);
fulladd full56 (sum[326], carry[326], 1'b0, 1'b0, 1'b0);
fulladd full57 (sum[327], carry[327], 1'b0, 1'b0, 1'b0);
fulladd full58 (sum[328], carry[328], 1'b0, 1'b0, 1'b0);
fulladd full59 (sum[329], carry[329], 1'b0, 1'b0, 1'b0);
fulladd full510 (sum[330], carry[330], 1'b0, 1'b0, 1'b0);
fulladd full511 (sum[331], carry[331], 1'b0, 1'b0, 1'b0);
fulladd full512 (sum[332], carry[332], 1'b0, 1'b0, 1'b0);
fulladd full513 (sum[333], carry[333], 1'b0, 1'b0, 1'b0);
fulladd full514 (sum[334], carry[334], 1'b0, 1'b0, 1'b0);
fulladd full515 (sum[335], carry[335], C[480], 1'b0, 1'b0);
fulladd full516 (sum[336], carry[336], C[481], C[512], 1'b0);
fulladd full517 (sum[337], carry[337], C[482], C[513], C[544]);
fulladd full518 (sum[338], carry[338], C[483], C[514], C[545]);
fulladd full519 (sum[339], carry[339], C[484], C[515], C[546]);
fulladd full520 (sum[340], carry[340], C[485], C[516], C[547]);
fulladd full521 (sum[341], carry[341], C[486], C[517], C[548]);
fulladd full522 (sum[342], carry[342], C[487], C[518], C[549]);
fulladd full523 (sum[343], carry[343], C[488], C[519], C[550]);
fulladd full524 (sum[344], carry[344], C[489], C[520], C[551]);
fulladd full525 (sum[345], carry[345], C[490], C[521], C[552]);
fulladd full526 (sum[346], carry[346], C[491], C[522], C[553]);
fulladd full527 (sum[347], carry[347], C[492], C[523], C[554]);
fulladd full528 (sum[348], carry[348], C[493], C[524], C[555]);
fulladd full529 (sum[349], carry[349], C[494], C[525], C[556]);
fulladd full530 (sum[350], carry[350], C[495], C[526], C[557]);
fulladd full531 (sum[351], carry[351], C[496], C[527], C[558]);
fulladd full532 (sum[352], carry[352], C[497], C[528], C[559]);
fulladd full533 (sum[353], carry[353], C[498], C[529], C[560]);
fulladd full534 (sum[354], carry[354], C[499], C[530], C[561]);
fulladd full535 (sum[355], carry[355], C[500], C[531], C[562]);
fulladd full536 (sum[356], carry[356], C[501], C[532], C[563]);
fulladd full537 (sum[357], carry[357], C[502], C[533], C[564]);
fulladd full538 (sum[358], carry[358], C[503], C[534], C[565]);
fulladd full539 (sum[359], carry[359], C[504], C[535], C[566]);
fulladd full540 (sum[360], carry[360], C[505], C[536], C[567]);
fulladd full541 (sum[361], carry[361], C[506], C[537], C[568]);
fulladd full542 (sum[362], carry[362], C[507], C[538], C[569]);
fulladd full543 (sum[363], carry[363], C[508], C[539], C[570]);
fulladd full544 (sum[364], carry[364], C[509], C[540], C[571]);
fulladd full545 (sum[365], carry[365], C[510], C[541], C[572]);
fulladd full546 (sum[366], carry[366], C[511], C[542], C[573]);
fulladd full547 (sum[367], carry[367], 1'b0, C[543], C[574]);
fulladd full548 (sum[368], carry[368], 1'b0, 1'b0, C[575]);
fulladd full549 (sum[369], carry[369], 1'b0, 1'b0, 1'b0);
fulladd full550 (sum[370], carry[370], 1'b0, 1'b0, 1'b0);
fulladd full551 (sum[371], carry[371], 1'b0, 1'b0, 1'b0);
fulladd full552 (sum[372], carry[372], 1'b0, 1'b0, 1'b0);
fulladd full553 (sum[373], carry[373], 1'b0, 1'b0, 1'b0);
fulladd full554 (sum[374], carry[374], 1'b0, 1'b0, 1'b0);
fulladd full555 (sum[375], carry[375], 1'b0, 1'b0, 1'b0);
fulladd full556 (sum[376], carry[376], 1'b0, 1'b0, 1'b0);
fulladd full557 (sum[377], carry[377], 1'b0, 1'b0, 1'b0);
fulladd full558 (sum[378], carry[378], 1'b0, 1'b0, 1'b0);
fulladd full559 (sum[379], carry[379], 1'b0, 1'b0, 1'b0);
fulladd full560 (sum[380], carry[380], 1'b0, 1'b0, 1'b0);
fulladd full561 (sum[381], carry[381], 1'b0, 1'b0, 1'b0);
fulladd full562 (sum[382], carry[382], 1'b0, 1'b0, 1'b0);
fulladd full563 (sum[383], carry[383], 1'b0, 1'b0, 1'b0);

//pp18,19,20
fulladd full60 (sum[384], carry[384], 1'b0, 1'b0, 1'b0);
fulladd full61 (sum[385], carry[385], 1'b0, 1'b0, 1'b0);
fulladd full62 (sum[386], carry[386], 1'b0, 1'b0, 1'b0);
fulladd full63 (sum[387], carry[387], 1'b0, 1'b0, 1'b0);
fulladd full64 (sum[388], carry[388], 1'b0, 1'b0, 1'b0);
fulladd full65 (sum[389], carry[389], 1'b0, 1'b0, 1'b0);
fulladd full66 (sum[390], carry[390], 1'b0, 1'b0, 1'b0);
fulladd full67 (sum[391], carry[391], 1'b0, 1'b0, 1'b0);
fulladd full68 (sum[392], carry[392], 1'b0, 1'b0, 1'b0);
fulladd full69 (sum[393], carry[393], 1'b0, 1'b0, 1'b0);
fulladd full610 (sum[394], carry[394], 1'b0, 1'b0, 1'b0);
fulladd full611 (sum[395], carry[395], 1'b0, 1'b0, 1'b0);
fulladd full612 (sum[396], carry[396], 1'b0, 1'b0, 1'b0);
fulladd full613 (sum[397], carry[397], 1'b0, 1'b0, 1'b0);
fulladd full614 (sum[398], carry[398], 1'b0, 1'b0, 1'b0);
fulladd full615 (sum[399], carry[399], 1'b0, 1'b0, 1'b0);
fulladd full616 (sum[400], carry[400], 1'b0, 1'b0, 1'b0);
fulladd full617 (sum[401], carry[401], 1'b0, 1'b0, 1'b0);
fulladd full618 (sum[402], carry[402], C[576], 1'b0, 1'b0);
fulladd full619 (sum[403], carry[403], C[577], C[608], 1'b0);
fulladd full620 (sum[404], carry[404], C[578], C[609], C[640]);
fulladd full621 (sum[405], carry[405], C[579], C[610], C[641]);
fulladd full622 (sum[406], carry[406], C[580], C[611], C[642]);
fulladd full623 (sum[407], carry[407], C[581], C[612], C[643]);
fulladd full624 (sum[408], carry[408], C[582], C[613], C[644]);
fulladd full625 (sum[409], carry[409], C[583], C[614], C[645]);
fulladd full626 (sum[410], carry[410], C[584], C[615], C[646]);
fulladd full627 (sum[411], carry[411], C[585], C[616], C[647]);
fulladd full628 (sum[412], carry[412], C[586], C[617], C[648]);
fulladd full629 (sum[413], carry[413], C[587], C[618], C[649]);
fulladd full630 (sum[414], carry[414], C[588], C[619], C[650]);
fulladd full631 (sum[415], carry[415], C[589], C[620], C[651]);
fulladd full632 (sum[416], carry[416], C[590], C[621], C[652]);
fulladd full633 (sum[417], carry[417], C[591], C[622], C[653]);
fulladd full634 (sum[418], carry[418], C[592], C[623], C[654]);
fulladd full635 (sum[419], carry[419], C[593], C[624], C[655]);
fulladd full636 (sum[420], carry[420], C[594], C[625], C[656]);
fulladd full637 (sum[421], carry[421], C[595], C[626], C[657]);
fulladd full638 (sum[422], carry[422], C[596], C[627], C[658]);
fulladd full639 (sum[423], carry[423], C[597], C[628], C[659]);
fulladd full640 (sum[424], carry[424], C[598], C[629], C[660]);
fulladd full641 (sum[425], carry[425], C[599], C[630], C[661]);
fulladd full642 (sum[426], carry[426], C[600], C[631], C[662]);
fulladd full643 (sum[427], carry[427], C[601], C[632], C[663]);
fulladd full644 (sum[428], carry[428], C[602], C[633], C[664]);
fulladd full645 (sum[429], carry[429], C[603], C[634], C[665]);
fulladd full646 (sum[430], carry[430], C[604], C[635], C[666]);
fulladd full647 (sum[431], carry[431], C[605], C[636], C[667]);
fulladd full648 (sum[432], carry[432], C[606], C[637], C[668]);
fulladd full649 (sum[433], carry[433], 1'b0, C[638], C[669]);
fulladd full650 (sum[434], carry[434], 1'b0, 1'b0, C[670]);
fulladd full651 (sum[435], carry[435], 1'b0, 1'b0, 1'b0);
fulladd full652 (sum[436], carry[436], 1'b0, 1'b0, 1'b0);
fulladd full653 (sum[437], carry[437], 1'b0, 1'b0, 1'b0);
fulladd full654 (sum[438], carry[438], 1'b0, 1'b0, 1'b0);
fulladd full655 (sum[439], carry[439], 1'b0, 1'b0, 1'b0);
fulladd full656 (sum[440], carry[440], 1'b0, 1'b0, 1'b0);
fulladd full657 (sum[441], carry[441], 1'b0, 1'b0, 1'b0);
fulladd full658 (sum[442], carry[442], 1'b0, 1'b0, 1'b0);
fulladd full659 (sum[443], carry[443], 1'b0, 1'b0, 1'b0);
fulladd full660 (sum[444], carry[444], 1'b0, 1'b0, 1'b0);
fulladd full661 (sum[445], carry[445], 1'b0, 1'b0, 1'b0);
fulladd full662 (sum[446], carry[446], 1'b0, 1'b0, 1'b0);
fulladd full663 (sum[447], carry[447], 1'b0, 1'b0, 1'b0);

//pp21,22,23
fulladd full70 (sum[448], carry[448], 1'b0, 1'b0, 1'b0);
fulladd full71 (sum[449], carry[449], 1'b0, 1'b0, 1'b0);
fulladd full72 (sum[450], carry[450], 1'b0, 1'b0, 1'b0);
fulladd full73 (sum[451], carry[451], 1'b0, 1'b0, 1'b0);
fulladd full74 (sum[452], carry[452], 1'b0, 1'b0, 1'b0);
fulladd full75 (sum[453], carry[453], 1'b0, 1'b0, 1'b0);
fulladd full76 (sum[454], carry[454], 1'b0, 1'b0, 1'b0);
fulladd full77 (sum[455], carry[455], 1'b0, 1'b0, 1'b0);
fulladd full78 (sum[456], carry[456], 1'b0, 1'b0, 1'b0);
fulladd full79 (sum[457], carry[457], 1'b0, 1'b0, 1'b0);
fulladd full710 (sum[458], carry[458], 1'b0, 1'b0, 1'b0);
fulladd full711 (sum[459], carry[459], 1'b0, 1'b0, 1'b0);
fulladd full712 (sum[460], carry[460], 1'b0, 1'b0, 1'b0);
fulladd full713 (sum[461], carry[461], 1'b0, 1'b0, 1'b0);
fulladd full714 (sum[462], carry[462], 1'b0, 1'b0, 1'b0);
fulladd full715 (sum[463], carry[463], 1'b0, 1'b0, 1'b0);
fulladd full716 (sum[464], carry[464], 1'b0, 1'b0, 1'b0);
fulladd full717 (sum[465], carry[465], 1'b0, 1'b0, 1'b0);
fulladd full718 (sum[466], carry[466], 1'b0, 1'b0, 1'b0);
fulladd full719 (sum[467], carry[467], 1'b0, 1'b0, 1'b0);
fulladd full720 (sum[468], carry[468], 1'b0, 1'b0, 1'b0);
fulladd full721 (sum[469], carry[469], C[672], 1'b0, 1'b0);
fulladd full722 (sum[470], carry[470], C[673], C[704], 1'b0);
fulladd full723 (sum[471], carry[471], C[674], C[705], C[736]);
fulladd full724 (sum[472], carry[472], C[675], C[706], C[737]);
fulladd full725 (sum[473], carry[473], C[676], C[707], C[738]);
fulladd full726 (sum[474], carry[474], C[677], C[708], C[739]);
fulladd full727 (sum[475], carry[475], C[678], C[709], C[740]);
fulladd full728 (sum[476], carry[476], C[679], C[710], C[741]);
fulladd full729 (sum[477], carry[477], C[680], C[711], C[742]);
fulladd full730 (sum[478], carry[478], C[681], C[712], C[743]);
fulladd full731 (sum[479], carry[479], C[682], C[713], C[744]);
fulladd full732 (sum[480], carry[480], C[683], C[714], C[745]);
fulladd full733 (sum[481], carry[481], C[684], C[715], C[746]);
fulladd full734 (sum[482], carry[482], C[685], C[716], C[747]);
fulladd full735 (sum[483], carry[483], C[686], C[717], C[748]);
fulladd full736 (sum[484], carry[484], C[687], C[718], C[749]);
fulladd full737 (sum[485], carry[485], C[688], C[719], C[750]);
fulladd full738 (sum[486], carry[486], C[689], C[720], C[751]);
fulladd full739 (sum[487], carry[487], C[690], C[721], C[752]);
fulladd full740 (sum[488], carry[488], C[691], C[722], C[753]);
fulladd full741 (sum[489], carry[489], C[692], C[723], C[754]);
fulladd full742 (sum[490], carry[490], C[693], C[724], C[755]);
fulladd full743 (sum[491], carry[491], C[694], C[725], C[756]);
fulladd full744 (sum[492], carry[492], C[695], C[726], C[757]);
fulladd full745 (sum[493], carry[493], C[696], C[727], C[758]);
fulladd full746 (sum[494], carry[494], C[697], C[728], C[759]);
fulladd full747 (sum[495], carry[495], C[698], C[729], C[760]);
fulladd full748 (sum[496], carry[496], C[699], C[730], C[761]);
fulladd full749 (sum[497], carry[497], C[700], C[731], C[762]);
fulladd full750 (sum[498], carry[498], C[701], C[732], C[763]);
fulladd full751 (sum[499], carry[499], C[702], C[733], C[764]);
fulladd full752 (sum[500], carry[500], C[703], C[734], C[765]);
fulladd full753 (sum[501], carry[501], 1'b0, C[735], C[766]);
fulladd full754 (sum[502], carry[502], 1'b0, 1'b0, C[767]);
fulladd full755 (sum[503], carry[503], 1'b0, 1'b0, 1'b0);
fulladd full756 (sum[504], carry[504], 1'b0, 1'b0, 1'b0);
fulladd full757 (sum[505], carry[505], 1'b0, 1'b0, 1'b0);
fulladd full758 (sum[506], carry[506], 1'b0, 1'b0, 1'b0);
fulladd full759 (sum[507], carry[507], 1'b0, 1'b0, 1'b0);
fulladd full760 (sum[508], carry[508], 1'b0, 1'b0, 1'b0);
fulladd full761 (sum[509], carry[509], 1'b0, 1'b0, 1'b0);
fulladd full762 (sum[510], carry[510], 1'b0, 1'b0, 1'b0);
fulladd full763 (sum[511], carry[511], 1'b0, 1'b0, 1'b0);

//pp24,25,26
fulladd full80 (sum[512], carry[512], 1'b0, 1'b0, 1'b0);
fulladd full81 (sum[513], carry[513], 1'b0, 1'b0, 1'b0);
fulladd full82 (sum[514], carry[514], 1'b0, 1'b0, 1'b0);
fulladd full83 (sum[515], carry[515], 1'b0, 1'b0, 1'b0);
fulladd full84 (sum[516], carry[516], 1'b0, 1'b0, 1'b0);
fulladd full85 (sum[517], carry[517], 1'b0, 1'b0, 1'b0);
fulladd full86 (sum[518], carry[518], 1'b0, 1'b0, 1'b0);
fulladd full87 (sum[519], carry[519], 1'b0, 1'b0, 1'b0);
fulladd full88 (sum[520], carry[520], 1'b0, 1'b0, 1'b0);
fulladd full89 (sum[521], carry[521], 1'b0, 1'b0, 1'b0);
fulladd full810 (sum[522], carry[522], 1'b0, 1'b0, 1'b0);
fulladd full811 (sum[523], carry[523], 1'b0, 1'b0, 1'b0);
fulladd full812 (sum[524], carry[524], 1'b0, 1'b0, 1'b0);
fulladd full813 (sum[525], carry[525], 1'b0, 1'b0, 1'b0);
fulladd full814 (sum[526], carry[526], 1'b0, 1'b0, 1'b0);
fulladd full815 (sum[527], carry[527], 1'b0, 1'b0, 1'b0);
fulladd full816 (sum[528], carry[528], 1'b0, 1'b0, 1'b0);
fulladd full817 (sum[529], carry[529], 1'b0, 1'b0, 1'b0);
fulladd full818 (sum[530], carry[530], 1'b0, 1'b0, 1'b0);
fulladd full819 (sum[531], carry[531], 1'b0, 1'b0, 1'b0);
fulladd full820 (sum[532], carry[532], 1'b0, 1'b0, 1'b0);
fulladd full821 (sum[533], carry[533], 1'b0, 1'b0, 1'b0);
fulladd full822 (sum[534], carry[534], 1'b0, 1'b0, 1'b0);
fulladd full823 (sum[535], carry[535], 1'b0, 1'b0, 1'b0);
fulladd full824 (sum[536], carry[536], C[768], 1'b0, 1'b0);
fulladd full825 (sum[537], carry[537], C[769], C[800], 1'b0);
fulladd full826 (sum[538], carry[538], C[770], C[801], C[832]);
fulladd full827 (sum[539], carry[539], C[771], C[802], C[833]);
fulladd full828 (sum[540], carry[540], C[772], C[803], C[834]);
fulladd full829 (sum[541], carry[541], C[773], C[804], C[835]);
fulladd full830 (sum[542], carry[542], C[774], C[805], C[836]);
fulladd full831 (sum[543], carry[543], C[775], C[806], C[837]);
fulladd full832 (sum[544], carry[544], C[776], C[807], C[838]);
fulladd full833 (sum[545], carry[545], C[777], C[808], C[839]);
fulladd full834 (sum[546], carry[546], C[778], C[809], C[840]);
fulladd full835 (sum[547], carry[547], C[779], C[810], C[841]);
fulladd full836 (sum[548], carry[548], C[780], C[811], C[842]);
fulladd full837 (sum[549], carry[549], C[781], C[812], C[843]);
fulladd full838 (sum[550], carry[550], C[782], C[813], C[844]);
fulladd full839 (sum[551], carry[551], C[783], C[814], C[845]);
fulladd full840 (sum[552], carry[552], C[784], C[815], C[846]);
fulladd full841 (sum[553], carry[553], C[785], C[816], C[847]);
fulladd full842 (sum[554], carry[554], C[786], C[817], C[848]);
fulladd full843 (sum[555], carry[555], C[787], C[818], C[849]);
fulladd full844 (sum[556], carry[556], C[788], C[819], C[850]);
fulladd full845 (sum[557], carry[557], C[789], C[820], C[851]);
fulladd full846 (sum[558], carry[558], C[790], C[821], C[852]);
fulladd full847 (sum[559], carry[559], C[791], C[822], C[853]);
fulladd full848 (sum[560], carry[560], C[792], C[823], C[854]);
fulladd full849 (sum[561], carry[561], C[793], C[824], C[855]);
fulladd full850 (sum[562], carry[562], C[794], C[825], C[856]);
fulladd full851 (sum[563], carry[563], C[795], C[826], C[857]);
fulladd full852 (sum[564], carry[564], C[796], C[827], C[858]);
fulladd full853 (sum[565], carry[565], C[797], C[828], C[859]);
fulladd full854 (sum[566], carry[566], C[798], C[829], C[860]);
fulladd full855 (sum[567], carry[567], C[799], C[830], C[861]);
fulladd full856 (sum[568], carry[568], 1'b0, C[831], C[862]);
fulladd full857 (sum[569], carry[569], 1'b0, 1'b0, C[863]);
fulladd full858 (sum[570], carry[570], 1'b0, 1'b0, 1'b0);
fulladd full859 (sum[571], carry[571], 1'b0, 1'b0, 1'b0);
fulladd full860 (sum[572], carry[572], 1'b0, 1'b0, 1'b0);
fulladd full861 (sum[573], carry[573], 1'b0, 1'b0, 1'b0);
fulladd full862 (sum[574], carry[574], 1'b0, 1'b0, 1'b0);
fulladd full863 (sum[575], carry[575], 1'b0, 1'b0, 1'b0);

//pp27,28,29
fulladd full90 (sum[576], carry[576], 1'b0, 1'b0, 1'b0);
fulladd full91 (sum[577], carry[577], 1'b0, 1'b0, 1'b0);
fulladd full92 (sum[578], carry[578], 1'b0, 1'b0, 1'b0);
fulladd full93 (sum[579], carry[579], 1'b0, 1'b0, 1'b0);
fulladd full94 (sum[580], carry[580], 1'b0, 1'b0, 1'b0);
fulladd full95 (sum[581], carry[581], 1'b0, 1'b0, 1'b0);
fulladd full96 (sum[582], carry[582], 1'b0, 1'b0, 1'b0);
fulladd full97 (sum[583], carry[583], 1'b0, 1'b0, 1'b0);
fulladd full98 (sum[584], carry[584], 1'b0, 1'b0, 1'b0);
fulladd full99 (sum[585], carry[585], 1'b0, 1'b0, 1'b0);
fulladd full910 (sum[586], carry[586], 1'b0, 1'b0, 1'b0);
fulladd full911 (sum[587], carry[587], 1'b0, 1'b0, 1'b0);
fulladd full912 (sum[588], carry[588], 1'b0, 1'b0, 1'b0);
fulladd full913 (sum[589], carry[589], 1'b0, 1'b0, 1'b0);
fulladd full914 (sum[590], carry[590], 1'b0, 1'b0, 1'b0);
fulladd full915 (sum[591], carry[591], 1'b0, 1'b0, 1'b0);
fulladd full916 (sum[592], carry[592], 1'b0, 1'b0, 1'b0);
fulladd full917 (sum[593], carry[593], 1'b0, 1'b0, 1'b0);
fulladd full918 (sum[594], carry[594], 1'b0, 1'b0, 1'b0);
fulladd full919 (sum[595], carry[595], 1'b0, 1'b0, 1'b0);
fulladd full920 (sum[596], carry[596], 1'b0, 1'b0, 1'b0);
fulladd full921 (sum[597], carry[597], 1'b0, 1'b0, 1'b0);
fulladd full922 (sum[598], carry[598], 1'b0, 1'b0, 1'b0);
fulladd full923 (sum[599], carry[599], 1'b0, 1'b0, 1'b0);
fulladd full924 (sum[600], carry[600], 1'b0, 1'b0, 1'b0);
fulladd full925 (sum[601], carry[601], 1'b0, 1'b0, 1'b0);
fulladd full926 (sum[602], carry[602], 1'b0, 1'b0, 1'b0);
fulladd full927 (sum[603], carry[603], C[864], 1'b0, 1'b0);
fulladd full928 (sum[604], carry[604], C[865], C[896], 1'b0);
fulladd full929 (sum[605], carry[605], C[866], C[897], C[928]);
fulladd full930 (sum[606], carry[606], C[867], C[898], C[929]);
fulladd full931 (sum[607], carry[607], C[868], C[899], C[930]);
fulladd full932 (sum[608], carry[608], C[869], C[900], C[931]);
fulladd full933 (sum[609], carry[609], C[870], C[901], C[932]);
fulladd full934 (sum[610], carry[610], C[871], C[902], C[933]);
fulladd full935 (sum[611], carry[611], C[872], C[903], C[934]);
fulladd full936 (sum[612], carry[612], C[873], C[904], C[935]);
fulladd full937 (sum[613], carry[613], C[874], C[905], C[936]);
fulladd full938 (sum[614], carry[614], C[875], C[906], C[937]);
fulladd full939 (sum[615], carry[615], C[876], C[907], C[938]);
fulladd full940 (sum[616], carry[616], C[877], C[908], C[939]);
fulladd full941 (sum[617], carry[617], C[878], C[909], C[940]);
fulladd full942 (sum[618], carry[618], C[879], C[910], C[941]);
fulladd full943 (sum[619], carry[619], C[880], C[911], C[942]);
fulladd full944 (sum[620], carry[620], C[881], C[912], C[943]);
fulladd full945 (sum[621], carry[621], C[882], C[913], C[944]);
fulladd full946 (sum[622], carry[622], C[883], C[914], C[945]);
fulladd full947 (sum[623], carry[623], C[884], C[915], C[946]);
fulladd full948 (sum[624], carry[624], C[885], C[916], C[947]);
fulladd full949 (sum[625], carry[625], C[886], C[917], C[948]);
fulladd full950 (sum[626], carry[626], C[887], C[918], C[949]);
fulladd full951 (sum[627], carry[627], C[888], C[919], C[950]);
fulladd full952 (sum[628], carry[628], C[889], C[920], C[951]);
fulladd full953 (sum[629], carry[629], C[890], C[921], C[952]);
fulladd full954 (sum[630], carry[630], C[891], C[922], C[953]);
fulladd full955 (sum[631], carry[631], C[892], C[923], C[954]);
fulladd full956 (sum[632], carry[632], C[893], C[924], C[955]);
fulladd full957 (sum[633], carry[633], C[894], C[925], C[956]);
fulladd full958 (sum[634], carry[634], C[895], C[926], C[957]);
fulladd full959 (sum[635], carry[635], 1'b0, C[927], C[958]);
fulladd full960 (sum[636], carry[636], 1'b0, 1'b0, C[959]);
fulladd full961 (sum[637], carry[637], 1'b0, 1'b0, 1'b0);
fulladd full962 (sum[638], carry[638], 1'b0, 1'b0, 1'b0);
fulladd full963 (sum[639], carry[639], 1'b0, 1'b0, 1'b0);

//sum0/1/2
fulladd full1_00 (sum_1[0], carry_1[0], sum[0], sum[64], sum[128]);
fulladd full1_01 (sum_1[1], carry_1[1], sum[1], sum[65], sum[129]);
fulladd full1_02 (sum_1[2], carry_1[2], sum[2], sum[66], sum[130]);
fulladd full1_03 (sum_1[3], carry_1[3], sum[3], sum[67], sum[131]);
fulladd full1_04 (sum_1[4], carry_1[4], sum[4], sum[68], sum[132]);
fulladd full1_05 (sum_1[5], carry_1[5], sum[5], sum[69], sum[133]);
fulladd full1_06 (sum_1[6], carry_1[6], sum[6], sum[70], sum[134]);
fulladd full1_07 (sum_1[7], carry_1[7], sum[7], sum[71], sum[135]);
fulladd full1_08 (sum_1[8], carry_1[8], sum[8], sum[72], sum[136]);
fulladd full1_09 (sum_1[9], carry_1[9], sum[9], sum[73], sum[137]);
fulladd full1_010 (sum_1[10], carry_1[10], sum[10], sum[74], sum[138]);
fulladd full1_011 (sum_1[11], carry_1[11], sum[11], sum[75], sum[139]);
fulladd full1_012 (sum_1[12], carry_1[12], sum[12], sum[76], sum[140]);
fulladd full1_013 (sum_1[13], carry_1[13], sum[13], sum[77], sum[141]);
fulladd full1_014 (sum_1[14], carry_1[14], sum[14], sum[78], sum[142]);
fulladd full1_015 (sum_1[15], carry_1[15], sum[15], sum[79], sum[143]);
fulladd full1_016 (sum_1[16], carry_1[16], sum[16], sum[80], sum[144]);
fulladd full1_017 (sum_1[17], carry_1[17], sum[17], sum[81], sum[145]);
fulladd full1_018 (sum_1[18], carry_1[18], sum[18], sum[82], sum[146]);
fulladd full1_019 (sum_1[19], carry_1[19], sum[19], sum[83], sum[147]);
fulladd full1_020 (sum_1[20], carry_1[20], sum[20], sum[84], sum[148]);
fulladd full1_021 (sum_1[21], carry_1[21], sum[21], sum[85], sum[149]);
fulladd full1_022 (sum_1[22], carry_1[22], sum[22], sum[86], sum[150]);
fulladd full1_023 (sum_1[23], carry_1[23], sum[23], sum[87], sum[151]);
fulladd full1_024 (sum_1[24], carry_1[24], sum[24], sum[88], sum[152]);
fulladd full1_025 (sum_1[25], carry_1[25], sum[25], sum[89], sum[153]);
fulladd full1_026 (sum_1[26], carry_1[26], sum[26], sum[90], sum[154]);
fulladd full1_027 (sum_1[27], carry_1[27], sum[27], sum[91], sum[155]);
fulladd full1_028 (sum_1[28], carry_1[28], sum[28], sum[92], sum[156]);
fulladd full1_029 (sum_1[29], carry_1[29], sum[29], sum[93], sum[157]);
fulladd full1_030 (sum_1[30], carry_1[30], sum[30], sum[94], sum[158]);
fulladd full1_031 (sum_1[31], carry_1[31], sum[31], sum[95], sum[159]);
fulladd full1_032 (sum_1[32], carry_1[32], sum[32], sum[96], sum[160]);
fulladd full1_033 (sum_1[33], carry_1[33], sum[33], sum[97], sum[161]);
fulladd full1_034 (sum_1[34], carry_1[34], sum[34], sum[98], sum[162]);
fulladd full1_035 (sum_1[35], carry_1[35], sum[35], sum[99], sum[163]);
fulladd full1_036 (sum_1[36], carry_1[36], sum[36], sum[100], sum[164]);
fulladd full1_037 (sum_1[37], carry_1[37], sum[37], sum[101], sum[165]);
fulladd full1_038 (sum_1[38], carry_1[38], sum[38], sum[102], sum[166]);
fulladd full1_039 (sum_1[39], carry_1[39], sum[39], sum[103], sum[167]);
fulladd full1_040 (sum_1[40], carry_1[40], sum[40], sum[104], sum[168]);
fulladd full1_041 (sum_1[41], carry_1[41], sum[41], sum[105], sum[169]);
fulladd full1_042 (sum_1[42], carry_1[42], sum[42], sum[106], sum[170]);
fulladd full1_043 (sum_1[43], carry_1[43], sum[43], sum[107], sum[171]);
fulladd full1_044 (sum_1[44], carry_1[44], sum[44], sum[108], sum[172]);
fulladd full1_045 (sum_1[45], carry_1[45], sum[45], sum[109], sum[173]);
fulladd full1_046 (sum_1[46], carry_1[46], sum[46], sum[110], sum[174]);
fulladd full1_047 (sum_1[47], carry_1[47], sum[47], sum[111], sum[175]);
fulladd full1_048 (sum_1[48], carry_1[48], sum[48], sum[112], sum[176]);
fulladd full1_049 (sum_1[49], carry_1[49], sum[49], sum[113], sum[177]);
fulladd full1_050 (sum_1[50], carry_1[50], sum[50], sum[114], sum[178]);
fulladd full1_051 (sum_1[51], carry_1[51], sum[51], sum[115], sum[179]);
fulladd full1_052 (sum_1[52], carry_1[52], sum[52], sum[116], sum[180]);
fulladd full1_053 (sum_1[53], carry_1[53], sum[53], sum[117], sum[181]);
fulladd full1_054 (sum_1[54], carry_1[54], sum[54], sum[118], sum[182]);
fulladd full1_055 (sum_1[55], carry_1[55], sum[55], sum[119], sum[183]);
fulladd full1_056 (sum_1[56], carry_1[56], sum[56], sum[120], sum[184]);
fulladd full1_057 (sum_1[57], carry_1[57], sum[57], sum[121], sum[185]);
fulladd full1_058 (sum_1[58], carry_1[58], sum[58], sum[122], sum[186]);
fulladd full1_059 (sum_1[59], carry_1[59], sum[59], sum[123], sum[187]);
fulladd full1_060 (sum_1[60], carry_1[60], sum[60], sum[124], sum[188]);
fulladd full1_061 (sum_1[61], carry_1[61], sum[61], sum[125], sum[189]);
fulladd full1_062 (sum_1[62], carry_1[62], sum[62], sum[126], sum[190]);
fulladd full1_063 (sum_1[63], carry_1[63], sum[63], sum[127], sum[191]);


//sum3/4/5
fulladd full1_10 (sum_1[64], carry_1[64], sum[192], sum[256], sum[320]);
fulladd full1_11 (sum_1[65], carry_1[65], sum[193], sum[257], sum[321]);
fulladd full1_12 (sum_1[66], carry_1[66], sum[194], sum[258], sum[322]);
fulladd full1_13 (sum_1[67], carry_1[67], sum[195], sum[259], sum[323]);
fulladd full1_14 (sum_1[68], carry_1[68], sum[196], sum[260], sum[324]);
fulladd full1_15 (sum_1[69], carry_1[69], sum[197], sum[261], sum[325]);
fulladd full1_16 (sum_1[70], carry_1[70], sum[198], sum[262], sum[326]);
fulladd full1_17 (sum_1[71], carry_1[71], sum[199], sum[263], sum[327]);
fulladd full1_18 (sum_1[72], carry_1[72], sum[200], sum[264], sum[328]);
fulladd full1_19 (sum_1[73], carry_1[73], sum[201], sum[265], sum[329]);
fulladd full1_110 (sum_1[74], carry_1[74], sum[202], sum[266], sum[330]);
fulladd full1_111 (sum_1[75], carry_1[75], sum[203], sum[267], sum[331]);
fulladd full1_112 (sum_1[76], carry_1[76], sum[204], sum[268], sum[332]);
fulladd full1_113 (sum_1[77], carry_1[77], sum[205], sum[269], sum[333]);
fulladd full1_114 (sum_1[78], carry_1[78], sum[206], sum[270], sum[334]);
fulladd full1_115 (sum_1[79], carry_1[79], sum[207], sum[271], sum[335]);
fulladd full1_116 (sum_1[80], carry_1[80], sum[208], sum[272], sum[336]);
fulladd full1_117 (sum_1[81], carry_1[81], sum[209], sum[273], sum[337]);
fulladd full1_118 (sum_1[82], carry_1[82], sum[210], sum[274], sum[338]);
fulladd full1_119 (sum_1[83], carry_1[83], sum[211], sum[275], sum[339]);
fulladd full1_120 (sum_1[84], carry_1[84], sum[212], sum[276], sum[340]);
fulladd full1_121 (sum_1[85], carry_1[85], sum[213], sum[277], sum[341]);
fulladd full1_122 (sum_1[86], carry_1[86], sum[214], sum[278], sum[342]);
fulladd full1_123 (sum_1[87], carry_1[87], sum[215], sum[279], sum[343]);
fulladd full1_124 (sum_1[88], carry_1[88], sum[216], sum[280], sum[344]);
fulladd full1_125 (sum_1[89], carry_1[89], sum[217], sum[281], sum[345]);
fulladd full1_126 (sum_1[90], carry_1[90], sum[218], sum[282], sum[346]);
fulladd full1_127 (sum_1[91], carry_1[91], sum[219], sum[283], sum[347]);
fulladd full1_128 (sum_1[92], carry_1[92], sum[220], sum[284], sum[348]);
fulladd full1_129 (sum_1[93], carry_1[93], sum[221], sum[285], sum[349]);
fulladd full1_130 (sum_1[94], carry_1[94], sum[222], sum[286], sum[350]);
fulladd full1_131 (sum_1[95], carry_1[95], sum[223], sum[287], sum[351]);
fulladd full1_132 (sum_1[96], carry_1[96], sum[224], sum[288], sum[352]);
fulladd full1_133 (sum_1[97], carry_1[97], sum[225], sum[289], sum[353]);
fulladd full1_134 (sum_1[98], carry_1[98], sum[226], sum[290], sum[354]);
fulladd full1_135 (sum_1[99], carry_1[99], sum[227], sum[291], sum[355]);
fulladd full1_136 (sum_1[100], carry_1[100], sum[228], sum[292], sum[356]);
fulladd full1_137 (sum_1[101], carry_1[101], sum[229], sum[293], sum[357]);
fulladd full1_138 (sum_1[102], carry_1[102], sum[230], sum[294], sum[358]);
fulladd full1_139 (sum_1[103], carry_1[103], sum[231], sum[295], sum[359]);
fulladd full1_140 (sum_1[104], carry_1[104], sum[232], sum[296], sum[360]);
fulladd full1_141 (sum_1[105], carry_1[105], sum[233], sum[297], sum[361]);
fulladd full1_142 (sum_1[106], carry_1[106], sum[234], sum[298], sum[362]);
fulladd full1_143 (sum_1[107], carry_1[107], sum[235], sum[299], sum[363]);
fulladd full1_144 (sum_1[108], carry_1[108], sum[236], sum[300], sum[364]);
fulladd full1_145 (sum_1[109], carry_1[109], sum[237], sum[301], sum[365]);
fulladd full1_146 (sum_1[110], carry_1[110], sum[238], sum[302], sum[366]);
fulladd full1_147 (sum_1[111], carry_1[111], sum[239], sum[303], sum[367]);
fulladd full1_148 (sum_1[112], carry_1[112], sum[240], sum[304], sum[368]);
fulladd full1_149 (sum_1[113], carry_1[113], sum[241], sum[305], sum[369]);
fulladd full1_150 (sum_1[114], carry_1[114], sum[242], sum[306], sum[370]);
fulladd full1_151 (sum_1[115], carry_1[115], sum[243], sum[307], sum[371]);
fulladd full1_152 (sum_1[116], carry_1[116], sum[244], sum[308], sum[372]);
fulladd full1_153 (sum_1[117], carry_1[117], sum[245], sum[309], sum[373]);
fulladd full1_154 (sum_1[118], carry_1[118], sum[246], sum[310], sum[374]);
fulladd full1_155 (sum_1[119], carry_1[119], sum[247], sum[311], sum[375]);
fulladd full1_156 (sum_1[120], carry_1[120], sum[248], sum[312], sum[376]);
fulladd full1_157 (sum_1[121], carry_1[121], sum[249], sum[313], sum[377]);
fulladd full1_158 (sum_1[122], carry_1[122], sum[250], sum[314], sum[378]);
fulladd full1_159 (sum_1[123], carry_1[123], sum[251], sum[315], sum[379]);
fulladd full1_160 (sum_1[124], carry_1[124], sum[252], sum[316], sum[380]);
fulladd full1_161 (sum_1[125], carry_1[125], sum[253], sum[317], sum[381]);
fulladd full1_162 (sum_1[126], carry_1[126], sum[254], sum[318], sum[382]);
fulladd full1_163 (sum_1[127], carry_1[127], sum[255], sum[319], sum[383]);

//sum6/7/8
fulladd full1_20 (sum_1[128], carry_1[128], sum[384], sum[448], sum[512]);
fulladd full1_21 (sum_1[129], carry_1[129], sum[385], sum[449], sum[513]);
fulladd full1_22 (sum_1[130], carry_1[130], sum[386], sum[450], sum[514]);
fulladd full1_23 (sum_1[131], carry_1[131], sum[387], sum[451], sum[515]);
fulladd full1_24 (sum_1[132], carry_1[132], sum[388], sum[452], sum[516]);
fulladd full1_25 (sum_1[133], carry_1[133], sum[389], sum[453], sum[517]);
fulladd full1_26 (sum_1[134], carry_1[134], sum[390], sum[454], sum[518]);
fulladd full1_27 (sum_1[135], carry_1[135], sum[391], sum[455], sum[519]);
fulladd full1_28 (sum_1[136], carry_1[136], sum[392], sum[456], sum[520]);
fulladd full1_29 (sum_1[137], carry_1[137], sum[393], sum[457], sum[521]);
fulladd full1_210 (sum_1[138], carry_1[138], sum[394], sum[458], sum[522]);
fulladd full1_211 (sum_1[139], carry_1[139], sum[395], sum[459], sum[523]);
fulladd full1_212 (sum_1[140], carry_1[140], sum[396], sum[460], sum[524]);
fulladd full1_213 (sum_1[141], carry_1[141], sum[397], sum[461], sum[525]);
fulladd full1_214 (sum_1[142], carry_1[142], sum[398], sum[462], sum[526]);
fulladd full1_215 (sum_1[143], carry_1[143], sum[399], sum[463], sum[527]);
fulladd full1_216 (sum_1[144], carry_1[144], sum[400], sum[464], sum[528]);
fulladd full1_217 (sum_1[145], carry_1[145], sum[401], sum[465], sum[529]);
fulladd full1_218 (sum_1[146], carry_1[146], sum[402], sum[466], sum[530]);
fulladd full1_219 (sum_1[147], carry_1[147], sum[403], sum[467], sum[531]);
fulladd full1_220 (sum_1[148], carry_1[148], sum[404], sum[468], sum[532]);
fulladd full1_221 (sum_1[149], carry_1[149], sum[405], sum[469], sum[533]);
fulladd full1_222 (sum_1[150], carry_1[150], sum[406], sum[470], sum[534]);
fulladd full1_223 (sum_1[151], carry_1[151], sum[407], sum[471], sum[535]);
fulladd full1_224 (sum_1[152], carry_1[152], sum[408], sum[472], sum[536]);
fulladd full1_225 (sum_1[153], carry_1[153], sum[409], sum[473], sum[537]);
fulladd full1_226 (sum_1[154], carry_1[154], sum[410], sum[474], sum[538]);
fulladd full1_227 (sum_1[155], carry_1[155], sum[411], sum[475], sum[539]);
fulladd full1_228 (sum_1[156], carry_1[156], sum[412], sum[476], sum[540]);
fulladd full1_229 (sum_1[157], carry_1[157], sum[413], sum[477], sum[541]);
fulladd full1_230 (sum_1[158], carry_1[158], sum[414], sum[478], sum[542]);
fulladd full1_231 (sum_1[159], carry_1[159], sum[415], sum[479], sum[543]);
fulladd full1_232 (sum_1[160], carry_1[160], sum[416], sum[480], sum[544]);
fulladd full1_233 (sum_1[161], carry_1[161], sum[417], sum[481], sum[545]);
fulladd full1_234 (sum_1[162], carry_1[162], sum[418], sum[482], sum[546]);
fulladd full1_235 (sum_1[163], carry_1[163], sum[419], sum[483], sum[547]);
fulladd full1_236 (sum_1[164], carry_1[164], sum[420], sum[484], sum[548]);
fulladd full1_237 (sum_1[165], carry_1[165], sum[421], sum[485], sum[549]);
fulladd full1_238 (sum_1[166], carry_1[166], sum[422], sum[486], sum[550]);
fulladd full1_239 (sum_1[167], carry_1[167], sum[423], sum[487], sum[551]);
fulladd full1_240 (sum_1[168], carry_1[168], sum[424], sum[488], sum[552]);
fulladd full1_241 (sum_1[169], carry_1[169], sum[425], sum[489], sum[553]);
fulladd full1_242 (sum_1[170], carry_1[170], sum[426], sum[490], sum[554]);
fulladd full1_243 (sum_1[171], carry_1[171], sum[427], sum[491], sum[555]);
fulladd full1_244 (sum_1[172], carry_1[172], sum[428], sum[492], sum[556]);
fulladd full1_245 (sum_1[173], carry_1[173], sum[429], sum[493], sum[557]);
fulladd full1_246 (sum_1[174], carry_1[174], sum[430], sum[494], sum[558]);
fulladd full1_247 (sum_1[175], carry_1[175], sum[431], sum[495], sum[559]);
fulladd full1_248 (sum_1[176], carry_1[176], sum[432], sum[496], sum[560]);
fulladd full1_249 (sum_1[177], carry_1[177], sum[433], sum[497], sum[561]);
fulladd full1_250 (sum_1[178], carry_1[178], sum[434], sum[498], sum[562]);
fulladd full1_251 (sum_1[179], carry_1[179], sum[435], sum[499], sum[563]);
fulladd full1_252 (sum_1[180], carry_1[180], sum[436], sum[500], sum[564]);
fulladd full1_253 (sum_1[181], carry_1[181], sum[437], sum[501], sum[565]);
fulladd full1_254 (sum_1[182], carry_1[182], sum[438], sum[502], sum[566]);
fulladd full1_255 (sum_1[183], carry_1[183], sum[439], sum[503], sum[567]);
fulladd full1_256 (sum_1[184], carry_1[184], sum[440], sum[504], sum[568]);
fulladd full1_257 (sum_1[185], carry_1[185], sum[441], sum[505], sum[569]);
fulladd full1_258 (sum_1[186], carry_1[186], sum[442], sum[506], sum[570]);
fulladd full1_259 (sum_1[187], carry_1[187], sum[443], sum[507], sum[571]);
fulladd full1_260 (sum_1[188], carry_1[188], sum[444], sum[508], sum[572]);
fulladd full1_261 (sum_1[189], carry_1[189], sum[445], sum[509], sum[573]);
fulladd full1_262 (sum_1[190], carry_1[190], sum[446], sum[510], sum[574]);
fulladd full1_263 (sum_1[191], carry_1[191], sum[447], sum[511], sum[575]);

//carry0/1/2
fulladd full1_30 (sum_1[192], carry_1[192], 1'b0, 1'b0, 1'b0);
fulladd full1_31 (sum_1[193], carry_1[193], carry[0], carry[64], carry[128]);
fulladd full1_32 (sum_1[194], carry_1[194], carry[1], carry[65], carry[129]);
fulladd full1_33 (sum_1[195], carry_1[195], carry[2], carry[66], carry[130]);
fulladd full1_34 (sum_1[196], carry_1[196], carry[3], carry[67], carry[131]);
fulladd full1_35 (sum_1[197], carry_1[197], carry[4], carry[68], carry[132]);
fulladd full1_36 (sum_1[198], carry_1[198], carry[5], carry[69], carry[133]);
fulladd full1_37 (sum_1[199], carry_1[199], carry[6], carry[70], carry[134]);
fulladd full1_38 (sum_1[200], carry_1[200], carry[7], carry[71], carry[135]);
fulladd full1_39 (sum_1[201], carry_1[201], carry[8], carry[72], carry[136]);
fulladd full1_310 (sum_1[202], carry_1[202], carry[9], carry[73], carry[137]);
fulladd full1_311 (sum_1[203], carry_1[203], carry[10], carry[74], carry[138]);
fulladd full1_312 (sum_1[204], carry_1[204], carry[11], carry[75], carry[139]);
fulladd full1_313 (sum_1[205], carry_1[205], carry[12], carry[76], carry[140]);
fulladd full1_314 (sum_1[206], carry_1[206], carry[13], carry[77], carry[141]);
fulladd full1_315 (sum_1[207], carry_1[207], carry[14], carry[78], carry[142]);
fulladd full1_316 (sum_1[208], carry_1[208], carry[15], carry[79], carry[143]);
fulladd full1_317 (sum_1[209], carry_1[209], carry[16], carry[80], carry[144]);
fulladd full1_318 (sum_1[210], carry_1[210], carry[17], carry[81], carry[145]);
fulladd full1_319 (sum_1[211], carry_1[211], carry[18], carry[82], carry[146]);
fulladd full1_320 (sum_1[212], carry_1[212], carry[19], carry[83], carry[147]);
fulladd full1_321 (sum_1[213], carry_1[213], carry[20], carry[84], carry[148]);
fulladd full1_322 (sum_1[214], carry_1[214], carry[21], carry[85], carry[149]);
fulladd full1_323 (sum_1[215], carry_1[215], carry[22], carry[86], carry[150]);
fulladd full1_324 (sum_1[216], carry_1[216], carry[23], carry[87], carry[151]);
fulladd full1_325 (sum_1[217], carry_1[217], carry[24], carry[88], carry[152]);
fulladd full1_326 (sum_1[218], carry_1[218], carry[25], carry[89], carry[153]);
fulladd full1_327 (sum_1[219], carry_1[219], carry[26], carry[90], carry[154]);
fulladd full1_328 (sum_1[220], carry_1[220], carry[27], carry[91], carry[155]);
fulladd full1_329 (sum_1[221], carry_1[221], carry[28], carry[92], carry[156]);
fulladd full1_330 (sum_1[222], carry_1[222], carry[29], carry[93], carry[157]);
fulladd full1_331 (sum_1[223], carry_1[223], carry[30], carry[94], carry[158]);
fulladd full1_332 (sum_1[224], carry_1[224], carry[31], carry[95], carry[159]);
fulladd full1_333 (sum_1[225], carry_1[225], carry[32], carry[96], carry[160]);
fulladd full1_334 (sum_1[226], carry_1[226], carry[33], carry[97], carry[161]);
fulladd full1_335 (sum_1[227], carry_1[227], carry[34], carry[98], carry[162]);
fulladd full1_336 (sum_1[228], carry_1[228], carry[35], carry[99], carry[163]);
fulladd full1_337 (sum_1[229], carry_1[229], carry[36], carry[100], carry[164]);
fulladd full1_338 (sum_1[230], carry_1[230], carry[37], carry[101], carry[165]);
fulladd full1_339 (sum_1[231], carry_1[231], carry[38], carry[102], carry[166]);
fulladd full1_340 (sum_1[232], carry_1[232], carry[39], carry[103], carry[167]);
fulladd full1_341 (sum_1[233], carry_1[233], carry[40], carry[104], carry[168]);
fulladd full1_342 (sum_1[234], carry_1[234], carry[41], carry[105], carry[169]);
fulladd full1_343 (sum_1[235], carry_1[235], carry[42], carry[106], carry[170]);
fulladd full1_344 (sum_1[236], carry_1[236], carry[43], carry[107], carry[171]);
fulladd full1_345 (sum_1[237], carry_1[237], carry[44], carry[108], carry[172]);
fulladd full1_346 (sum_1[238], carry_1[238], carry[45], carry[109], carry[173]);
fulladd full1_347 (sum_1[239], carry_1[239], carry[46], carry[110], carry[174]);
fulladd full1_348 (sum_1[240], carry_1[240], carry[47], carry[111], carry[175]);
fulladd full1_349 (sum_1[241], carry_1[241], carry[48], carry[112], carry[176]);
fulladd full1_350 (sum_1[242], carry_1[242], carry[49], carry[113], carry[177]);
fulladd full1_351 (sum_1[243], carry_1[243], carry[50], carry[114], carry[178]);
fulladd full1_352 (sum_1[244], carry_1[244], carry[51], carry[115], carry[179]);
fulladd full1_353 (sum_1[245], carry_1[245], carry[52], carry[116], carry[180]);
fulladd full1_354 (sum_1[246], carry_1[246], carry[53], carry[117], carry[181]);
fulladd full1_355 (sum_1[247], carry_1[247], carry[54], carry[118], carry[182]);
fulladd full1_356 (sum_1[248], carry_1[248], carry[55], carry[119], carry[183]);
fulladd full1_357 (sum_1[249], carry_1[249], carry[56], carry[120], carry[184]);
fulladd full1_358 (sum_1[250], carry_1[250], carry[57], carry[121], carry[185]);
fulladd full1_359 (sum_1[251], carry_1[251], carry[58], carry[122], carry[186]);
fulladd full1_360 (sum_1[252], carry_1[252], carry[59], carry[123], carry[187]);
fulladd full1_361 (sum_1[253], carry_1[253], carry[60], carry[124], carry[188]);
fulladd full1_362 (sum_1[254], carry_1[254], carry[61], carry[125], carry[189]);
fulladd full1_363 (sum_1[255], carry_1[255], carry[62], carry[126], carry[190]);


//carry3/4/5
fulladd full1_40 (sum_1[256], carry_1[256], 1'b0, 1'b0, 1'b0);
fulladd full1_41 (sum_1[257], carry_1[257], carry[192], carry[256], carry[320]);
fulladd full1_42 (sum_1[258], carry_1[258], carry[193], carry[257], carry[321]);
fulladd full1_43 (sum_1[259], carry_1[259], carry[194], carry[258], carry[322]);
fulladd full1_44 (sum_1[260], carry_1[260], carry[195], carry[259], carry[323]);
fulladd full1_45 (sum_1[261], carry_1[261], carry[196], carry[260], carry[324]);
fulladd full1_46 (sum_1[262], carry_1[262], carry[197], carry[261], carry[325]);
fulladd full1_47 (sum_1[263], carry_1[263], carry[198], carry[262], carry[326]);
fulladd full1_48 (sum_1[264], carry_1[264], carry[199], carry[263], carry[327]);
fulladd full1_49 (sum_1[265], carry_1[265], carry[200], carry[264], carry[328]);
fulladd full1_410 (sum_1[266], carry_1[266], carry[201], carry[265], carry[329]);
fulladd full1_411 (sum_1[267], carry_1[267], carry[202], carry[266], carry[330]);
fulladd full1_412 (sum_1[268], carry_1[268], carry[203], carry[267], carry[331]);
fulladd full1_413 (sum_1[269], carry_1[269], carry[204], carry[268], carry[332]);
fulladd full1_414 (sum_1[270], carry_1[270], carry[205], carry[269], carry[333]);
fulladd full1_415 (sum_1[271], carry_1[271], carry[206], carry[270], carry[334]);
fulladd full1_416 (sum_1[272], carry_1[272], carry[207], carry[271], carry[335]);
fulladd full1_417 (sum_1[273], carry_1[273], carry[208], carry[272], carry[336]);
fulladd full1_418 (sum_1[274], carry_1[274], carry[209], carry[273], carry[337]);
fulladd full1_419 (sum_1[275], carry_1[275], carry[210], carry[274], carry[338]);
fulladd full1_420 (sum_1[276], carry_1[276], carry[211], carry[275], carry[339]);
fulladd full1_421 (sum_1[277], carry_1[277], carry[212], carry[276], carry[340]);
fulladd full1_422 (sum_1[278], carry_1[278], carry[213], carry[277], carry[341]);
fulladd full1_423 (sum_1[279], carry_1[279], carry[214], carry[278], carry[342]);
fulladd full1_424 (sum_1[280], carry_1[280], carry[215], carry[279], carry[343]);
fulladd full1_425 (sum_1[281], carry_1[281], carry[216], carry[280], carry[344]);
fulladd full1_426 (sum_1[282], carry_1[282], carry[217], carry[281], carry[345]);
fulladd full1_427 (sum_1[283], carry_1[283], carry[218], carry[282], carry[346]);
fulladd full1_428 (sum_1[284], carry_1[284], carry[219], carry[283], carry[347]);
fulladd full1_429 (sum_1[285], carry_1[285], carry[220], carry[284], carry[348]);
fulladd full1_430 (sum_1[286], carry_1[286], carry[221], carry[285], carry[349]);
fulladd full1_431 (sum_1[287], carry_1[287], carry[222], carry[286], carry[350]);
fulladd full1_432 (sum_1[288], carry_1[288], carry[223], carry[287], carry[351]);
fulladd full1_433 (sum_1[289], carry_1[289], carry[224], carry[288], carry[352]);
fulladd full1_434 (sum_1[290], carry_1[290], carry[225], carry[289], carry[353]);
fulladd full1_435 (sum_1[291], carry_1[291], carry[226], carry[290], carry[354]);
fulladd full1_436 (sum_1[292], carry_1[292], carry[227], carry[291], carry[355]);
fulladd full1_437 (sum_1[293], carry_1[293], carry[228], carry[292], carry[356]);
fulladd full1_438 (sum_1[294], carry_1[294], carry[229], carry[293], carry[357]);
fulladd full1_439 (sum_1[295], carry_1[295], carry[230], carry[294], carry[358]);
fulladd full1_440 (sum_1[296], carry_1[296], carry[231], carry[295], carry[359]);
fulladd full1_441 (sum_1[297], carry_1[297], carry[232], carry[296], carry[360]);
fulladd full1_442 (sum_1[298], carry_1[298], carry[233], carry[297], carry[361]);
fulladd full1_443 (sum_1[299], carry_1[299], carry[234], carry[298], carry[362]);
fulladd full1_444 (sum_1[300], carry_1[300], carry[235], carry[299], carry[363]);
fulladd full1_445 (sum_1[301], carry_1[301], carry[236], carry[300], carry[364]);
fulladd full1_446 (sum_1[302], carry_1[302], carry[237], carry[301], carry[365]);
fulladd full1_447 (sum_1[303], carry_1[303], carry[238], carry[302], carry[366]);
fulladd full1_448 (sum_1[304], carry_1[304], carry[239], carry[303], carry[367]);
fulladd full1_449 (sum_1[305], carry_1[305], carry[240], carry[304], carry[368]);
fulladd full1_450 (sum_1[306], carry_1[306], carry[241], carry[305], carry[369]);
fulladd full1_451 (sum_1[307], carry_1[307], carry[242], carry[306], carry[370]);
fulladd full1_452 (sum_1[308], carry_1[308], carry[243], carry[307], carry[371]);
fulladd full1_453 (sum_1[309], carry_1[309], carry[244], carry[308], carry[372]);
fulladd full1_454 (sum_1[310], carry_1[310], carry[245], carry[309], carry[373]);
fulladd full1_455 (sum_1[311], carry_1[311], carry[246], carry[310], carry[374]);
fulladd full1_456 (sum_1[312], carry_1[312], carry[247], carry[311], carry[375]);
fulladd full1_457 (sum_1[313], carry_1[313], carry[248], carry[312], carry[376]);
fulladd full1_458 (sum_1[314], carry_1[314], carry[249], carry[313], carry[377]);
fulladd full1_459 (sum_1[315], carry_1[315], carry[250], carry[314], carry[378]);
fulladd full1_460 (sum_1[316], carry_1[316], carry[251], carry[315], carry[379]);
fulladd full1_461 (sum_1[317], carry_1[317], carry[252], carry[316], carry[380]);
fulladd full1_462 (sum_1[318], carry_1[318], carry[253], carry[317], carry[381]);
fulladd full1_463 (sum_1[319], carry_1[319], carry[254], carry[318], carry[382]);

//carry6/7/8/
fulladd full1_50 (sum_1[320], carry_1[320], 1'b0, 1'b0, 1'b0);
fulladd full1_51 (sum_1[321], carry_1[321], carry[384], carry[448], carry[512]);
fulladd full1_52 (sum_1[322], carry_1[322], carry[385], carry[449], carry[513]);
fulladd full1_53 (sum_1[323], carry_1[323], carry[386], carry[450], carry[514]);
fulladd full1_54 (sum_1[324], carry_1[324], carry[387], carry[451], carry[515]);
fulladd full1_55 (sum_1[325], carry_1[325], carry[388], carry[452], carry[516]);
fulladd full1_56 (sum_1[326], carry_1[326], carry[389], carry[453], carry[517]);
fulladd full1_57 (sum_1[327], carry_1[327], carry[390], carry[454], carry[518]);
fulladd full1_58 (sum_1[328], carry_1[328], carry[391], carry[455], carry[519]);
fulladd full1_59 (sum_1[329], carry_1[329], carry[392], carry[456], carry[520]);
fulladd full1_510 (sum_1[330], carry_1[330], carry[393], carry[457], carry[521]);
fulladd full1_511 (sum_1[331], carry_1[331], carry[394], carry[458], carry[522]);
fulladd full1_512 (sum_1[332], carry_1[332], carry[395], carry[459], carry[523]);
fulladd full1_513 (sum_1[333], carry_1[333], carry[396], carry[460], carry[524]);
fulladd full1_514 (sum_1[334], carry_1[334], carry[397], carry[461], carry[525]);
fulladd full1_515 (sum_1[335], carry_1[335], carry[398], carry[462], carry[526]);
fulladd full1_516 (sum_1[336], carry_1[336], carry[399], carry[463], carry[527]);
fulladd full1_517 (sum_1[337], carry_1[337], carry[400], carry[464], carry[528]);
fulladd full1_518 (sum_1[338], carry_1[338], carry[401], carry[465], carry[529]);
fulladd full1_519 (sum_1[339], carry_1[339], carry[402], carry[466], carry[530]);
fulladd full1_520 (sum_1[340], carry_1[340], carry[403], carry[467], carry[531]);
fulladd full1_521 (sum_1[341], carry_1[341], carry[404], carry[468], carry[532]);
fulladd full1_522 (sum_1[342], carry_1[342], carry[405], carry[469], carry[533]);
fulladd full1_523 (sum_1[343], carry_1[343], carry[406], carry[470], carry[534]);
fulladd full1_524 (sum_1[344], carry_1[344], carry[407], carry[471], carry[535]);
fulladd full1_525 (sum_1[345], carry_1[345], carry[408], carry[472], carry[536]);
fulladd full1_526 (sum_1[346], carry_1[346], carry[409], carry[473], carry[537]);
fulladd full1_527 (sum_1[347], carry_1[347], carry[410], carry[474], carry[538]);
fulladd full1_528 (sum_1[348], carry_1[348], carry[411], carry[475], carry[539]);
fulladd full1_529 (sum_1[349], carry_1[349], carry[412], carry[476], carry[540]);
fulladd full1_530 (sum_1[350], carry_1[350], carry[413], carry[477], carry[541]);
fulladd full1_531 (sum_1[351], carry_1[351], carry[414], carry[478], carry[542]);
fulladd full1_532 (sum_1[352], carry_1[352], carry[415], carry[479], carry[543]);
fulladd full1_533 (sum_1[353], carry_1[353], carry[416], carry[480], carry[544]);
fulladd full1_534 (sum_1[354], carry_1[354], carry[417], carry[481], carry[545]);
fulladd full1_535 (sum_1[355], carry_1[355], carry[418], carry[482], carry[546]);
fulladd full1_536 (sum_1[356], carry_1[356], carry[419], carry[483], carry[547]);
fulladd full1_537 (sum_1[357], carry_1[357], carry[420], carry[484], carry[548]);
fulladd full1_538 (sum_1[358], carry_1[358], carry[421], carry[485], carry[549]);
fulladd full1_539 (sum_1[359], carry_1[359], carry[422], carry[486], carry[550]);
fulladd full1_540 (sum_1[360], carry_1[360], carry[423], carry[487], carry[551]);
fulladd full1_541 (sum_1[361], carry_1[361], carry[424], carry[488], carry[552]);
fulladd full1_542 (sum_1[362], carry_1[362], carry[425], carry[489], carry[553]);
fulladd full1_543 (sum_1[363], carry_1[363], carry[426], carry[490], carry[554]);
fulladd full1_544 (sum_1[364], carry_1[364], carry[427], carry[491], carry[555]);
fulladd full1_545 (sum_1[365], carry_1[365], carry[428], carry[492], carry[556]);
fulladd full1_546 (sum_1[366], carry_1[366], carry[429], carry[493], carry[557]);
fulladd full1_547 (sum_1[367], carry_1[367], carry[430], carry[494], carry[558]);
fulladd full1_548 (sum_1[368], carry_1[368], carry[431], carry[495], carry[559]);
fulladd full1_549 (sum_1[369], carry_1[369], carry[432], carry[496], carry[560]);
fulladd full1_550 (sum_1[370], carry_1[370], carry[433], carry[497], carry[561]);
fulladd full1_551 (sum_1[371], carry_1[371], carry[434], carry[498], carry[562]);
fulladd full1_552 (sum_1[372], carry_1[372], carry[435], carry[499], carry[563]);
fulladd full1_553 (sum_1[373], carry_1[373], carry[436], carry[500], carry[564]);
fulladd full1_554 (sum_1[374], carry_1[374], carry[437], carry[501], carry[565]);
fulladd full1_555 (sum_1[375], carry_1[375], carry[438], carry[502], carry[566]);
fulladd full1_556 (sum_1[376], carry_1[376], carry[439], carry[503], carry[567]);
fulladd full1_557 (sum_1[377], carry_1[377], carry[440], carry[504], carry[568]);
fulladd full1_558 (sum_1[378], carry_1[378], carry[441], carry[505], carry[569]);
fulladd full1_559 (sum_1[379], carry_1[379], carry[442], carry[506], carry[570]);
fulladd full1_560 (sum_1[380], carry_1[380], carry[443], carry[507], carry[571]);
fulladd full1_561 (sum_1[381], carry_1[381], carry[444], carry[508], carry[572]);
fulladd full1_562 (sum_1[382], carry_1[382], carry[445], carry[509], carry[573]);
fulladd full1_563 (sum_1[383], carry_1[383], carry[446], carry[510], carry[574]);


//sum9/carry9/pp30
fulladd full1_60 (sum_1[384], carry_1[384], sum[576], 1'b0, 1'b0);
fulladd full1_61 (sum_1[385], carry_1[385], sum[577], carry[576], 1'b0);
fulladd full1_62 (sum_1[386], carry_1[386], sum[578], carry[577], 1'b0);
fulladd full1_63 (sum_1[387], carry_1[387], sum[579], carry[578], 1'b0);
fulladd full1_64 (sum_1[388], carry_1[388], sum[580], carry[579], 1'b0);
fulladd full1_65 (sum_1[389], carry_1[389], sum[581], carry[580], 1'b0);
fulladd full1_66 (sum_1[390], carry_1[390], sum[582], carry[581], 1'b0);
fulladd full1_67 (sum_1[391], carry_1[391], sum[583], carry[582], 1'b0);
fulladd full1_68 (sum_1[392], carry_1[392], sum[584], carry[583], 1'b0);
fulladd full1_69 (sum_1[393], carry_1[393], sum[585], carry[584], 1'b0);
fulladd full1_610 (sum_1[394], carry_1[394], sum[586], carry[585], 1'b0);
fulladd full1_611 (sum_1[395], carry_1[395], sum[587], carry[586], 1'b0);
fulladd full1_612 (sum_1[396], carry_1[396], sum[588], carry[587], 1'b0);
fulladd full1_613 (sum_1[397], carry_1[397], sum[589], carry[588], 1'b0);
fulladd full1_614 (sum_1[398], carry_1[398], sum[590], carry[589], 1'b0);
fulladd full1_615 (sum_1[399], carry_1[399], sum[591], carry[590], 1'b0);
fulladd full1_616 (sum_1[400], carry_1[400], sum[592], carry[591], 1'b0);
fulladd full1_617 (sum_1[401], carry_1[401], sum[593], carry[592], 1'b0);
fulladd full1_618 (sum_1[402], carry_1[402], sum[594], carry[593], 1'b0);
fulladd full1_619 (sum_1[403], carry_1[403], sum[595], carry[594], 1'b0);
fulladd full1_620 (sum_1[404], carry_1[404], sum[596], carry[595], 1'b0);
fulladd full1_621 (sum_1[405], carry_1[405], sum[597], carry[596], 1'b0);
fulladd full1_622 (sum_1[406], carry_1[406], sum[598], carry[597], 1'b0);
fulladd full1_623 (sum_1[407], carry_1[407], sum[599], carry[598], 1'b0);
fulladd full1_624 (sum_1[408], carry_1[408], sum[600], carry[599], 1'b0);
fulladd full1_625 (sum_1[409], carry_1[409], sum[601], carry[600], 1'b0);
fulladd full1_626 (sum_1[410], carry_1[410], sum[602], carry[601], 1'b0);
fulladd full1_627 (sum_1[411], carry_1[411], sum[603], carry[602], 1'b0);
fulladd full1_628 (sum_1[412], carry_1[412], sum[604], carry[603], 1'b0);
fulladd full1_629 (sum_1[413], carry_1[413], sum[605], carry[604], 1'b0);
fulladd full1_630 (sum_1[414], carry_1[414], sum[606], carry[605], C[960]);
fulladd full1_631 (sum_1[415], carry_1[415], sum[607], carry[606], C[961]);
fulladd full1_632 (sum_1[416], carry_1[416], sum[608], carry[607], C[962]);
fulladd full1_633 (sum_1[417], carry_1[417], sum[609], carry[608], C[963]);
fulladd full1_634 (sum_1[418], carry_1[418], sum[610], carry[609], C[964]);
fulladd full1_635 (sum_1[419], carry_1[419], sum[611], carry[610], C[965]);
fulladd full1_636 (sum_1[420], carry_1[420], sum[612], carry[611], C[966]);
fulladd full1_637 (sum_1[421], carry_1[421], sum[613], carry[612], C[967]);
fulladd full1_638 (sum_1[422], carry_1[422], sum[614], carry[613], C[968]);
fulladd full1_639 (sum_1[423], carry_1[423], sum[615], carry[614], C[969]);
fulladd full1_640 (sum_1[424], carry_1[424], sum[616], carry[615], C[970]);
fulladd full1_641 (sum_1[425], carry_1[425], sum[617], carry[616], C[971]);
fulladd full1_642 (sum_1[426], carry_1[426], sum[618], carry[617], C[972]);
fulladd full1_643 (sum_1[427], carry_1[427], sum[619], carry[618], C[973]);
fulladd full1_644 (sum_1[428], carry_1[428], sum[620], carry[619], C[974]);
fulladd full1_645 (sum_1[429], carry_1[429], sum[621], carry[620], C[975]);
fulladd full1_646 (sum_1[430], carry_1[430], sum[622], carry[621], C[976]);
fulladd full1_647 (sum_1[431], carry_1[431], sum[623], carry[622], C[977]);
fulladd full1_648 (sum_1[432], carry_1[432], sum[624], carry[623], C[978]);
fulladd full1_649 (sum_1[433], carry_1[433], sum[625], carry[624], C[979]);
fulladd full1_650 (sum_1[434], carry_1[434], sum[626], carry[625], C[980]);
fulladd full1_651 (sum_1[435], carry_1[435], sum[627], carry[626], C[981]);
fulladd full1_652 (sum_1[436], carry_1[436], sum[628], carry[627], C[982]);
fulladd full1_653 (sum_1[437], carry_1[437], sum[629], carry[628], C[983]);
fulladd full1_654 (sum_1[438], carry_1[438], sum[630], carry[629], C[984]);
fulladd full1_655 (sum_1[439], carry_1[439], sum[631], carry[630], C[985]);
fulladd full1_656 (sum_1[440], carry_1[440], sum[632], carry[631], C[986]);
fulladd full1_657 (sum_1[441], carry_1[441], sum[633], carry[632], C[987]);
fulladd full1_658 (sum_1[442], carry_1[442], sum[634], carry[633], C[988]);
fulladd full1_659 (sum_1[443], carry_1[443], sum[635], carry[634], C[989]);
fulladd full1_660 (sum_1[444], carry_1[444], sum[636], carry[635], C[990]);
fulladd full1_661 (sum_1[445], carry_1[445], sum[637], carry[636], C[991]);
fulladd full1_662 (sum_1[446], carry_1[446], sum[638], carry[637], C[991]);
fulladd full1_663 (sum_1[447], carry_1[447], sum[639], carry[638], C[991]);

//sum_1/0/1/2
fulladd full2_00 (sum_2[0], carry_2[0], sum_1[0], sum_1[64], sum_1[128]);
fulladd full2_01 (sum_2[1], carry_2[1], sum_1[1], sum_1[65], sum_1[129]);
fulladd full2_02 (sum_2[2], carry_2[2], sum_1[2], sum_1[66], sum_1[130]);
fulladd full2_03 (sum_2[3], carry_2[3], sum_1[3], sum_1[67], sum_1[131]);
fulladd full2_04 (sum_2[4], carry_2[4], sum_1[4], sum_1[68], sum_1[132]);
fulladd full2_05 (sum_2[5], carry_2[5], sum_1[5], sum_1[69], sum_1[133]);
fulladd full2_06 (sum_2[6], carry_2[6], sum_1[6], sum_1[70], sum_1[134]);
fulladd full2_07 (sum_2[7], carry_2[7], sum_1[7], sum_1[71], sum_1[135]);
fulladd full2_08 (sum_2[8], carry_2[8], sum_1[8], sum_1[72], sum_1[136]);
fulladd full2_09 (sum_2[9], carry_2[9], sum_1[9], sum_1[73], sum_1[137]);
fulladd full2_010 (sum_2[10], carry_2[10], sum_1[10], sum_1[74], sum_1[138]);
fulladd full2_011 (sum_2[11], carry_2[11], sum_1[11], sum_1[75], sum_1[139]);
fulladd full2_012 (sum_2[12], carry_2[12], sum_1[12], sum_1[76], sum_1[140]);
fulladd full2_013 (sum_2[13], carry_2[13], sum_1[13], sum_1[77], sum_1[141]);
fulladd full2_014 (sum_2[14], carry_2[14], sum_1[14], sum_1[78], sum_1[142]);
fulladd full2_015 (sum_2[15], carry_2[15], sum_1[15], sum_1[79], sum_1[143]);
fulladd full2_016 (sum_2[16], carry_2[16], sum_1[16], sum_1[80], sum_1[144]);
fulladd full2_017 (sum_2[17], carry_2[17], sum_1[17], sum_1[81], sum_1[145]);
fulladd full2_018 (sum_2[18], carry_2[18], sum_1[18], sum_1[82], sum_1[146]);
fulladd full2_019 (sum_2[19], carry_2[19], sum_1[19], sum_1[83], sum_1[147]);
fulladd full2_020 (sum_2[20], carry_2[20], sum_1[20], sum_1[84], sum_1[148]);
fulladd full2_021 (sum_2[21], carry_2[21], sum_1[21], sum_1[85], sum_1[149]);
fulladd full2_022 (sum_2[22], carry_2[22], sum_1[22], sum_1[86], sum_1[150]);
fulladd full2_023 (sum_2[23], carry_2[23], sum_1[23], sum_1[87], sum_1[151]);
fulladd full2_024 (sum_2[24], carry_2[24], sum_1[24], sum_1[88], sum_1[152]);
fulladd full2_025 (sum_2[25], carry_2[25], sum_1[25], sum_1[89], sum_1[153]);
fulladd full2_026 (sum_2[26], carry_2[26], sum_1[26], sum_1[90], sum_1[154]);
fulladd full2_027 (sum_2[27], carry_2[27], sum_1[27], sum_1[91], sum_1[155]);
fulladd full2_028 (sum_2[28], carry_2[28], sum_1[28], sum_1[92], sum_1[156]);
fulladd full2_029 (sum_2[29], carry_2[29], sum_1[29], sum_1[93], sum_1[157]);
fulladd full2_030 (sum_2[30], carry_2[30], sum_1[30], sum_1[94], sum_1[158]);
fulladd full2_031 (sum_2[31], carry_2[31], sum_1[31], sum_1[95], sum_1[159]);
fulladd full2_032 (sum_2[32], carry_2[32], sum_1[32], sum_1[96], sum_1[160]);
fulladd full2_033 (sum_2[33], carry_2[33], sum_1[33], sum_1[97], sum_1[161]);
fulladd full2_034 (sum_2[34], carry_2[34], sum_1[34], sum_1[98], sum_1[162]);
fulladd full2_035 (sum_2[35], carry_2[35], sum_1[35], sum_1[99], sum_1[163]);
fulladd full2_036 (sum_2[36], carry_2[36], sum_1[36], sum_1[100], sum_1[164]);
fulladd full2_037 (sum_2[37], carry_2[37], sum_1[37], sum_1[101], sum_1[165]);
fulladd full2_038 (sum_2[38], carry_2[38], sum_1[38], sum_1[102], sum_1[166]);
fulladd full2_039 (sum_2[39], carry_2[39], sum_1[39], sum_1[103], sum_1[167]);
fulladd full2_040 (sum_2[40], carry_2[40], sum_1[40], sum_1[104], sum_1[168]);
fulladd full2_041 (sum_2[41], carry_2[41], sum_1[41], sum_1[105], sum_1[169]);
fulladd full2_042 (sum_2[42], carry_2[42], sum_1[42], sum_1[106], sum_1[170]);
fulladd full2_043 (sum_2[43], carry_2[43], sum_1[43], sum_1[107], sum_1[171]);
fulladd full2_044 (sum_2[44], carry_2[44], sum_1[44], sum_1[108], sum_1[172]);
fulladd full2_045 (sum_2[45], carry_2[45], sum_1[45], sum_1[109], sum_1[173]);
fulladd full2_046 (sum_2[46], carry_2[46], sum_1[46], sum_1[110], sum_1[174]);
fulladd full2_047 (sum_2[47], carry_2[47], sum_1[47], sum_1[111], sum_1[175]);
fulladd full2_048 (sum_2[48], carry_2[48], sum_1[48], sum_1[112], sum_1[176]);
fulladd full2_049 (sum_2[49], carry_2[49], sum_1[49], sum_1[113], sum_1[177]);
fulladd full2_050 (sum_2[50], carry_2[50], sum_1[50], sum_1[114], sum_1[178]);
fulladd full2_051 (sum_2[51], carry_2[51], sum_1[51], sum_1[115], sum_1[179]);
fulladd full2_052 (sum_2[52], carry_2[52], sum_1[52], sum_1[116], sum_1[180]);
fulladd full2_053 (sum_2[53], carry_2[53], sum_1[53], sum_1[117], sum_1[181]);
fulladd full2_054 (sum_2[54], carry_2[54], sum_1[54], sum_1[118], sum_1[182]);
fulladd full2_055 (sum_2[55], carry_2[55], sum_1[55], sum_1[119], sum_1[183]);
fulladd full2_056 (sum_2[56], carry_2[56], sum_1[56], sum_1[120], sum_1[184]);
fulladd full2_057 (sum_2[57], carry_2[57], sum_1[57], sum_1[121], sum_1[185]);
fulladd full2_058 (sum_2[58], carry_2[58], sum_1[58], sum_1[122], sum_1[186]);
fulladd full2_059 (sum_2[59], carry_2[59], sum_1[59], sum_1[123], sum_1[187]);
fulladd full2_060 (sum_2[60], carry_2[60], sum_1[60], sum_1[124], sum_1[188]);
fulladd full2_061 (sum_2[61], carry_2[61], sum_1[61], sum_1[125], sum_1[189]);
fulladd full2_062 (sum_2[62], carry_2[62], sum_1[62], sum_1[126], sum_1[190]);
fulladd full2_063 (sum_2[63], carry_2[63], sum_1[63], sum_1[127], sum_1[191]);

//sum_1/3/4/5
fulladd full2_10 (sum_2[64], carry_2[64], sum_1[192], sum_1[256], sum_1[320]);
fulladd full2_11 (sum_2[65], carry_2[65], sum_1[193], sum_1[257], sum_1[321]);
fulladd full2_12 (sum_2[66], carry_2[66], sum_1[194], sum_1[258], sum_1[322]);
fulladd full2_13 (sum_2[67], carry_2[67], sum_1[195], sum_1[259], sum_1[323]);
fulladd full2_14 (sum_2[68], carry_2[68], sum_1[196], sum_1[260], sum_1[324]);
fulladd full2_15 (sum_2[69], carry_2[69], sum_1[197], sum_1[261], sum_1[325]);
fulladd full2_16 (sum_2[70], carry_2[70], sum_1[198], sum_1[262], sum_1[326]);
fulladd full2_17 (sum_2[71], carry_2[71], sum_1[199], sum_1[263], sum_1[327]);
fulladd full2_18 (sum_2[72], carry_2[72], sum_1[200], sum_1[264], sum_1[328]);
fulladd full2_19 (sum_2[73], carry_2[73], sum_1[201], sum_1[265], sum_1[329]);
fulladd full2_110 (sum_2[74], carry_2[74], sum_1[202], sum_1[266], sum_1[330]);
fulladd full2_111 (sum_2[75], carry_2[75], sum_1[203], sum_1[267], sum_1[331]);
fulladd full2_112 (sum_2[76], carry_2[76], sum_1[204], sum_1[268], sum_1[332]);
fulladd full2_113 (sum_2[77], carry_2[77], sum_1[205], sum_1[269], sum_1[333]);
fulladd full2_114 (sum_2[78], carry_2[78], sum_1[206], sum_1[270], sum_1[334]);
fulladd full2_115 (sum_2[79], carry_2[79], sum_1[207], sum_1[271], sum_1[335]);
fulladd full2_116 (sum_2[80], carry_2[80], sum_1[208], sum_1[272], sum_1[336]);
fulladd full2_117 (sum_2[81], carry_2[81], sum_1[209], sum_1[273], sum_1[337]);
fulladd full2_118 (sum_2[82], carry_2[82], sum_1[210], sum_1[274], sum_1[338]);
fulladd full2_119 (sum_2[83], carry_2[83], sum_1[211], sum_1[275], sum_1[339]);
fulladd full2_120 (sum_2[84], carry_2[84], sum_1[212], sum_1[276], sum_1[340]);
fulladd full2_121 (sum_2[85], carry_2[85], sum_1[213], sum_1[277], sum_1[341]);
fulladd full2_122 (sum_2[86], carry_2[86], sum_1[214], sum_1[278], sum_1[342]);
fulladd full2_123 (sum_2[87], carry_2[87], sum_1[215], sum_1[279], sum_1[343]);
fulladd full2_124 (sum_2[88], carry_2[88], sum_1[216], sum_1[280], sum_1[344]);
fulladd full2_125 (sum_2[89], carry_2[89], sum_1[217], sum_1[281], sum_1[345]);
fulladd full2_126 (sum_2[90], carry_2[90], sum_1[218], sum_1[282], sum_1[346]);
fulladd full2_127 (sum_2[91], carry_2[91], sum_1[219], sum_1[283], sum_1[347]);
fulladd full2_128 (sum_2[92], carry_2[92], sum_1[220], sum_1[284], sum_1[348]);
fulladd full2_129 (sum_2[93], carry_2[93], sum_1[221], sum_1[285], sum_1[349]);
fulladd full2_130 (sum_2[94], carry_2[94], sum_1[222], sum_1[286], sum_1[350]);
fulladd full2_131 (sum_2[95], carry_2[95], sum_1[223], sum_1[287], sum_1[351]);
fulladd full2_132 (sum_2[96], carry_2[96], sum_1[224], sum_1[288], sum_1[352]);
fulladd full2_133 (sum_2[97], carry_2[97], sum_1[225], sum_1[289], sum_1[353]);
fulladd full2_134 (sum_2[98], carry_2[98], sum_1[226], sum_1[290], sum_1[354]);
fulladd full2_135 (sum_2[99], carry_2[99], sum_1[227], sum_1[291], sum_1[355]);
fulladd full2_136 (sum_2[100], carry_2[100], sum_1[228], sum_1[292], sum_1[356]);
fulladd full2_137 (sum_2[101], carry_2[101], sum_1[229], sum_1[293], sum_1[357]);
fulladd full2_138 (sum_2[102], carry_2[102], sum_1[230], sum_1[294], sum_1[358]);
fulladd full2_139 (sum_2[103], carry_2[103], sum_1[231], sum_1[295], sum_1[359]);
fulladd full2_140 (sum_2[104], carry_2[104], sum_1[232], sum_1[296], sum_1[360]);
fulladd full2_141 (sum_2[105], carry_2[105], sum_1[233], sum_1[297], sum_1[361]);
fulladd full2_142 (sum_2[106], carry_2[106], sum_1[234], sum_1[298], sum_1[362]);
fulladd full2_143 (sum_2[107], carry_2[107], sum_1[235], sum_1[299], sum_1[363]);
fulladd full2_144 (sum_2[108], carry_2[108], sum_1[236], sum_1[300], sum_1[364]);
fulladd full2_145 (sum_2[109], carry_2[109], sum_1[237], sum_1[301], sum_1[365]);
fulladd full2_146 (sum_2[110], carry_2[110], sum_1[238], sum_1[302], sum_1[366]);
fulladd full2_147 (sum_2[111], carry_2[111], sum_1[239], sum_1[303], sum_1[367]);
fulladd full2_148 (sum_2[112], carry_2[112], sum_1[240], sum_1[304], sum_1[368]);
fulladd full2_149 (sum_2[113], carry_2[113], sum_1[241], sum_1[305], sum_1[369]);
fulladd full2_150 (sum_2[114], carry_2[114], sum_1[242], sum_1[306], sum_1[370]);
fulladd full2_151 (sum_2[115], carry_2[115], sum_1[243], sum_1[307], sum_1[371]);
fulladd full2_152 (sum_2[116], carry_2[116], sum_1[244], sum_1[308], sum_1[372]);
fulladd full2_153 (sum_2[117], carry_2[117], sum_1[245], sum_1[309], sum_1[373]);
fulladd full2_154 (sum_2[118], carry_2[118], sum_1[246], sum_1[310], sum_1[374]);
fulladd full2_155 (sum_2[119], carry_2[119], sum_1[247], sum_1[311], sum_1[375]);
fulladd full2_156 (sum_2[120], carry_2[120], sum_1[248], sum_1[312], sum_1[376]);
fulladd full2_157 (sum_2[121], carry_2[121], sum_1[249], sum_1[313], sum_1[377]);
fulladd full2_158 (sum_2[122], carry_2[122], sum_1[250], sum_1[314], sum_1[378]);
fulladd full2_159 (sum_2[123], carry_2[123], sum_1[251], sum_1[315], sum_1[379]);
fulladd full2_160 (sum_2[124], carry_2[124], sum_1[252], sum_1[316], sum_1[380]);
fulladd full2_161 (sum_2[125], carry_2[125], sum_1[253], sum_1[317], sum_1[381]);
fulladd full2_162 (sum_2[126], carry_2[126], sum_1[254], sum_1[318], sum_1[382]);
fulladd full2_163 (sum_2[127], carry_2[127], sum_1[255], sum_1[319], sum_1[383]);

//carry_1/0/1/2
fulladd full2_20 (sum_2[128], carry_2[128], 1'b0, 1'b0, 1'b0);
fulladd full2_21 (sum_2[129], carry_2[129], carry_1[0], carry_1[64], carry_1[128]);
fulladd full2_22 (sum_2[130], carry_2[130], carry_1[1], carry_1[65], carry_1[129]);
fulladd full2_23 (sum_2[131], carry_2[131], carry_1[2], carry_1[66], carry_1[130]);
fulladd full2_24 (sum_2[132], carry_2[132], carry_1[3], carry_1[67], carry_1[131]);
fulladd full2_25 (sum_2[133], carry_2[133], carry_1[4], carry_1[68], carry_1[132]);
fulladd full2_26 (sum_2[134], carry_2[134], carry_1[5], carry_1[69], carry_1[133]);
fulladd full2_27 (sum_2[135], carry_2[135], carry_1[6], carry_1[70], carry_1[134]);
fulladd full2_28 (sum_2[136], carry_2[136], carry_1[7], carry_1[71], carry_1[135]);
fulladd full2_29 (sum_2[137], carry_2[137], carry_1[8], carry_1[72], carry_1[136]);
fulladd full2_210 (sum_2[138], carry_2[138], carry_1[9], carry_1[73], carry_1[137]);
fulladd full2_211 (sum_2[139], carry_2[139], carry_1[10], carry_1[74], carry_1[138]);
fulladd full2_212 (sum_2[140], carry_2[140], carry_1[11], carry_1[75], carry_1[139]);
fulladd full2_213 (sum_2[141], carry_2[141], carry_1[12], carry_1[76], carry_1[140]);
fulladd full2_214 (sum_2[142], carry_2[142], carry_1[13], carry_1[77], carry_1[141]);
fulladd full2_215 (sum_2[143], carry_2[143], carry_1[14], carry_1[78], carry_1[142]);
fulladd full2_216 (sum_2[144], carry_2[144], carry_1[15], carry_1[79], carry_1[143]);
fulladd full2_217 (sum_2[145], carry_2[145], carry_1[16], carry_1[80], carry_1[144]);
fulladd full2_218 (sum_2[146], carry_2[146], carry_1[17], carry_1[81], carry_1[145]);
fulladd full2_219 (sum_2[147], carry_2[147], carry_1[18], carry_1[82], carry_1[146]);
fulladd full2_220 (sum_2[148], carry_2[148], carry_1[19], carry_1[83], carry_1[147]);
fulladd full2_221 (sum_2[149], carry_2[149], carry_1[20], carry_1[84], carry_1[148]);
fulladd full2_222 (sum_2[150], carry_2[150], carry_1[21], carry_1[85], carry_1[149]);
fulladd full2_223 (sum_2[151], carry_2[151], carry_1[22], carry_1[86], carry_1[150]);
fulladd full2_224 (sum_2[152], carry_2[152], carry_1[23], carry_1[87], carry_1[151]);
fulladd full2_225 (sum_2[153], carry_2[153], carry_1[24], carry_1[88], carry_1[152]);
fulladd full2_226 (sum_2[154], carry_2[154], carry_1[25], carry_1[89], carry_1[153]);
fulladd full2_227 (sum_2[155], carry_2[155], carry_1[26], carry_1[90], carry_1[154]);
fulladd full2_228 (sum_2[156], carry_2[156], carry_1[27], carry_1[91], carry_1[155]);
fulladd full2_229 (sum_2[157], carry_2[157], carry_1[28], carry_1[92], carry_1[156]);
fulladd full2_230 (sum_2[158], carry_2[158], carry_1[29], carry_1[93], carry_1[157]);
fulladd full2_231 (sum_2[159], carry_2[159], carry_1[30], carry_1[94], carry_1[158]);
fulladd full2_232 (sum_2[160], carry_2[160], carry_1[31], carry_1[95], carry_1[159]);
fulladd full2_233 (sum_2[161], carry_2[161], carry_1[32], carry_1[96], carry_1[160]);
fulladd full2_234 (sum_2[162], carry_2[162], carry_1[33], carry_1[97], carry_1[161]);
fulladd full2_235 (sum_2[163], carry_2[163], carry_1[34], carry_1[98], carry_1[162]);
fulladd full2_236 (sum_2[164], carry_2[164], carry_1[35], carry_1[99], carry_1[163]);
fulladd full2_237 (sum_2[165], carry_2[165], carry_1[36], carry_1[100], carry_1[164]);
fulladd full2_238 (sum_2[166], carry_2[166], carry_1[37], carry_1[101], carry_1[165]);
fulladd full2_239 (sum_2[167], carry_2[167], carry_1[38], carry_1[102], carry_1[166]);
fulladd full2_240 (sum_2[168], carry_2[168], carry_1[39], carry_1[103], carry_1[167]);
fulladd full2_241 (sum_2[169], carry_2[169], carry_1[40], carry_1[104], carry_1[168]);
fulladd full2_242 (sum_2[170], carry_2[170], carry_1[41], carry_1[105], carry_1[169]);
fulladd full2_243 (sum_2[171], carry_2[171], carry_1[42], carry_1[106], carry_1[170]);
fulladd full2_244 (sum_2[172], carry_2[172], carry_1[43], carry_1[107], carry_1[171]);
fulladd full2_245 (sum_2[173], carry_2[173], carry_1[44], carry_1[108], carry_1[172]);
fulladd full2_246 (sum_2[174], carry_2[174], carry_1[45], carry_1[109], carry_1[173]);
fulladd full2_247 (sum_2[175], carry_2[175], carry_1[46], carry_1[110], carry_1[174]);
fulladd full2_248 (sum_2[176], carry_2[176], carry_1[47], carry_1[111], carry_1[175]);
fulladd full2_249 (sum_2[177], carry_2[177], carry_1[48], carry_1[112], carry_1[176]);
fulladd full2_250 (sum_2[178], carry_2[178], carry_1[49], carry_1[113], carry_1[177]);
fulladd full2_251 (sum_2[179], carry_2[179], carry_1[50], carry_1[114], carry_1[178]);
fulladd full2_252 (sum_2[180], carry_2[180], carry_1[51], carry_1[115], carry_1[179]);
fulladd full2_253 (sum_2[181], carry_2[181], carry_1[52], carry_1[116], carry_1[180]);
fulladd full2_254 (sum_2[182], carry_2[182], carry_1[53], carry_1[117], carry_1[181]);
fulladd full2_255 (sum_2[183], carry_2[183], carry_1[54], carry_1[118], carry_1[182]);
fulladd full2_256 (sum_2[184], carry_2[184], carry_1[55], carry_1[119], carry_1[183]);
fulladd full2_257 (sum_2[185], carry_2[185], carry_1[56], carry_1[120], carry_1[184]);
fulladd full2_258 (sum_2[186], carry_2[186], carry_1[57], carry_1[121], carry_1[185]);
fulladd full2_259 (sum_2[187], carry_2[187], carry_1[58], carry_1[122], carry_1[186]);
fulladd full2_260 (sum_2[188], carry_2[188], carry_1[59], carry_1[123], carry_1[187]);
fulladd full2_261 (sum_2[189], carry_2[189], carry_1[60], carry_1[124], carry_1[188]);
fulladd full2_262 (sum_2[190], carry_2[190], carry_1[61], carry_1[125], carry_1[189]);
fulladd full2_263 (sum_2[191], carry_2[191], carry_1[62], carry_1[126], carry_1[190]);

//carry_1/3/4/5
fulladd full2_30 (sum_2[192], carry_2[192], 1'b0, 1'b0, 1'b0);
fulladd full2_31 (sum_2[193], carry_2[193], carry_1[192], carry_1[256], carry_1[320]);
fulladd full2_32 (sum_2[194], carry_2[194], carry_1[193], carry_1[257], carry_1[321]);
fulladd full2_33 (sum_2[195], carry_2[195], carry_1[194], carry_1[258], carry_1[322]);
fulladd full2_34 (sum_2[196], carry_2[196], carry_1[195], carry_1[259], carry_1[323]);
fulladd full2_35 (sum_2[197], carry_2[197], carry_1[196], carry_1[260], carry_1[324]);
fulladd full2_36 (sum_2[198], carry_2[198], carry_1[197], carry_1[261], carry_1[325]);
fulladd full2_37 (sum_2[199], carry_2[199], carry_1[198], carry_1[262], carry_1[326]);
fulladd full2_38 (sum_2[200], carry_2[200], carry_1[199], carry_1[263], carry_1[327]);
fulladd full2_39 (sum_2[201], carry_2[201], carry_1[200], carry_1[264], carry_1[328]);
fulladd full2_310 (sum_2[202], carry_2[202], carry_1[201], carry_1[265], carry_1[329]);
fulladd full2_311 (sum_2[203], carry_2[203], carry_1[202], carry_1[266], carry_1[330]);
fulladd full2_312 (sum_2[204], carry_2[204], carry_1[203], carry_1[267], carry_1[331]);
fulladd full2_313 (sum_2[205], carry_2[205], carry_1[204], carry_1[268], carry_1[332]);
fulladd full2_314 (sum_2[206], carry_2[206], carry_1[205], carry_1[269], carry_1[333]);
fulladd full2_315 (sum_2[207], carry_2[207], carry_1[206], carry_1[270], carry_1[334]);
fulladd full2_316 (sum_2[208], carry_2[208], carry_1[207], carry_1[271], carry_1[335]);
fulladd full2_317 (sum_2[209], carry_2[209], carry_1[208], carry_1[272], carry_1[336]);
fulladd full2_318 (sum_2[210], carry_2[210], carry_1[209], carry_1[273], carry_1[337]);
fulladd full2_319 (sum_2[211], carry_2[211], carry_1[210], carry_1[274], carry_1[338]);
fulladd full2_320 (sum_2[212], carry_2[212], carry_1[211], carry_1[275], carry_1[339]);
fulladd full2_321 (sum_2[213], carry_2[213], carry_1[212], carry_1[276], carry_1[340]);
fulladd full2_322 (sum_2[214], carry_2[214], carry_1[213], carry_1[277], carry_1[341]);
fulladd full2_323 (sum_2[215], carry_2[215], carry_1[214], carry_1[278], carry_1[342]);
fulladd full2_324 (sum_2[216], carry_2[216], carry_1[215], carry_1[279], carry_1[343]);
fulladd full2_325 (sum_2[217], carry_2[217], carry_1[216], carry_1[280], carry_1[344]);
fulladd full2_326 (sum_2[218], carry_2[218], carry_1[217], carry_1[281], carry_1[345]);
fulladd full2_327 (sum_2[219], carry_2[219], carry_1[218], carry_1[282], carry_1[346]);
fulladd full2_328 (sum_2[220], carry_2[220], carry_1[219], carry_1[283], carry_1[347]);
fulladd full2_329 (sum_2[221], carry_2[221], carry_1[220], carry_1[284], carry_1[348]);
fulladd full2_330 (sum_2[222], carry_2[222], carry_1[221], carry_1[285], carry_1[349]);
fulladd full2_331 (sum_2[223], carry_2[223], carry_1[222], carry_1[286], carry_1[350]);
fulladd full2_332 (sum_2[224], carry_2[224], carry_1[223], carry_1[287], carry_1[351]);
fulladd full2_333 (sum_2[225], carry_2[225], carry_1[224], carry_1[288], carry_1[352]);
fulladd full2_334 (sum_2[226], carry_2[226], carry_1[225], carry_1[289], carry_1[353]);
fulladd full2_335 (sum_2[227], carry_2[227], carry_1[226], carry_1[290], carry_1[354]);
fulladd full2_336 (sum_2[228], carry_2[228], carry_1[227], carry_1[291], carry_1[355]);
fulladd full2_337 (sum_2[229], carry_2[229], carry_1[228], carry_1[292], carry_1[356]);
fulladd full2_338 (sum_2[230], carry_2[230], carry_1[229], carry_1[293], carry_1[357]);
fulladd full2_339 (sum_2[231], carry_2[231], carry_1[230], carry_1[294], carry_1[358]);
fulladd full2_340 (sum_2[232], carry_2[232], carry_1[231], carry_1[295], carry_1[359]);
fulladd full2_341 (sum_2[233], carry_2[233], carry_1[232], carry_1[296], carry_1[360]);
fulladd full2_342 (sum_2[234], carry_2[234], carry_1[233], carry_1[297], carry_1[361]);
fulladd full2_343 (sum_2[235], carry_2[235], carry_1[234], carry_1[298], carry_1[362]);
fulladd full2_344 (sum_2[236], carry_2[236], carry_1[235], carry_1[299], carry_1[363]);
fulladd full2_345 (sum_2[237], carry_2[237], carry_1[236], carry_1[300], carry_1[364]);
fulladd full2_346 (sum_2[238], carry_2[238], carry_1[237], carry_1[301], carry_1[365]);
fulladd full2_347 (sum_2[239], carry_2[239], carry_1[238], carry_1[302], carry_1[366]);
fulladd full2_348 (sum_2[240], carry_2[240], carry_1[239], carry_1[303], carry_1[367]);
fulladd full2_349 (sum_2[241], carry_2[241], carry_1[240], carry_1[304], carry_1[368]);
fulladd full2_350 (sum_2[242], carry_2[242], carry_1[241], carry_1[305], carry_1[369]);
fulladd full2_351 (sum_2[243], carry_2[243], carry_1[242], carry_1[306], carry_1[370]);
fulladd full2_352 (sum_2[244], carry_2[244], carry_1[243], carry_1[307], carry_1[371]);
fulladd full2_353 (sum_2[245], carry_2[245], carry_1[244], carry_1[308], carry_1[372]);
fulladd full2_354 (sum_2[246], carry_2[246], carry_1[245], carry_1[309], carry_1[373]);
fulladd full2_355 (sum_2[247], carry_2[247], carry_1[246], carry_1[310], carry_1[374]);
fulladd full2_356 (sum_2[248], carry_2[248], carry_1[247], carry_1[311], carry_1[375]);
fulladd full2_357 (sum_2[249], carry_2[249], carry_1[248], carry_1[312], carry_1[376]);
fulladd full2_358 (sum_2[250], carry_2[250], carry_1[249], carry_1[313], carry_1[377]);
fulladd full2_359 (sum_2[251], carry_2[251], carry_1[250], carry_1[314], carry_1[378]);
fulladd full2_360 (sum_2[252], carry_2[252], carry_1[251], carry_1[315], carry_1[379]);
fulladd full2_361 (sum_2[253], carry_2[253], carry_1[252], carry_1[316], carry_1[380]);
fulladd full2_362 (sum_2[254], carry_2[254], carry_1[253], carry_1[317], carry_1[381]);
fulladd full2_363 (sum_2[255], carry_2[255], carry_1[254], carry_1[318], carry_1[382]);


//sum_1/6.carry_1/6.pp31
fulladd full2_40 (sum_2[256], carry_2[256], sum_1[384], 1'b0, 1'b0);
fulladd full2_41 (sum_2[257], carry_2[257], sum_1[385], carry_1[384], 1'b0);
fulladd full2_42 (sum_2[258], carry_2[258], sum_1[386], carry_1[385], 1'b0);
fulladd full2_43 (sum_2[259], carry_2[259], sum_1[387], carry_1[386], 1'b0);
fulladd full2_44 (sum_2[260], carry_2[260], sum_1[388], carry_1[387], 1'b0);
fulladd full2_45 (sum_2[261], carry_2[261], sum_1[389], carry_1[388], 1'b0);
fulladd full2_46 (sum_2[262], carry_2[262], sum_1[390], carry_1[389], 1'b0);
fulladd full2_47 (sum_2[263], carry_2[263], sum_1[391], carry_1[390], 1'b0);
fulladd full2_48 (sum_2[264], carry_2[264], sum_1[392], carry_1[391], 1'b0);
fulladd full2_49 (sum_2[265], carry_2[265], sum_1[393], carry_1[392], 1'b0);
fulladd full2_410 (sum_2[266], carry_2[266], sum_1[394], carry_1[393], 1'b0);
fulladd full2_411 (sum_2[267], carry_2[267], sum_1[395], carry_1[394], 1'b0);
fulladd full2_412 (sum_2[268], carry_2[268], sum_1[396], carry_1[395], 1'b0);
fulladd full2_413 (sum_2[269], carry_2[269], sum_1[397], carry_1[396], 1'b0);
fulladd full2_414 (sum_2[270], carry_2[270], sum_1[398], carry_1[397], 1'b0);
fulladd full2_415 (sum_2[271], carry_2[271], sum_1[399], carry_1[398], 1'b0);
fulladd full2_416 (sum_2[272], carry_2[272], sum_1[400], carry_1[399], 1'b0);
fulladd full2_417 (sum_2[273], carry_2[273], sum_1[401], carry_1[400], 1'b0);
fulladd full2_418 (sum_2[274], carry_2[274], sum_1[402], carry_1[401], 1'b0);
fulladd full2_419 (sum_2[275], carry_2[275], sum_1[403], carry_1[402], 1'b0);
fulladd full2_420 (sum_2[276], carry_2[276], sum_1[404], carry_1[403], 1'b0);
fulladd full2_421 (sum_2[277], carry_2[277], sum_1[405], carry_1[404], 1'b0);
fulladd full2_422 (sum_2[278], carry_2[278], sum_1[406], carry_1[405], 1'b0);
fulladd full2_423 (sum_2[279], carry_2[279], sum_1[407], carry_1[406], 1'b0);
fulladd full2_424 (sum_2[280], carry_2[280], sum_1[408], carry_1[407], 1'b0);
fulladd full2_425 (sum_2[281], carry_2[281], sum_1[409], carry_1[408], 1'b0);
fulladd full2_426 (sum_2[282], carry_2[282], sum_1[410], carry_1[409], 1'b0);
fulladd full2_427 (sum_2[283], carry_2[283], sum_1[411], carry_1[410], 1'b0);
fulladd full2_428 (sum_2[284], carry_2[284], sum_1[412], carry_1[411], 1'b0);
fulladd full2_429 (sum_2[285], carry_2[285], sum_1[413], carry_1[412], 1'b0);
fulladd full2_430 (sum_2[286], carry_2[286], sum_1[414], carry_1[413], 1'b0);
fulladd full2_431 (sum_2[287], carry_2[287], sum_1[415], carry_1[414], C[992]);
fulladd full2_432 (sum_2[288], carry_2[288], sum_1[416], carry_1[415], C[993]);
fulladd full2_433 (sum_2[289], carry_2[289], sum_1[417], carry_1[416], C[994]);
fulladd full2_434 (sum_2[290], carry_2[290], sum_1[418], carry_1[417], C[995]);
fulladd full2_435 (sum_2[291], carry_2[291], sum_1[419], carry_1[418], C[996]);
fulladd full2_436 (sum_2[292], carry_2[292], sum_1[420], carry_1[419], C[997]);
fulladd full2_437 (sum_2[293], carry_2[293], sum_1[421], carry_1[420], C[998]);
fulladd full2_438 (sum_2[294], carry_2[294], sum_1[422], carry_1[421], C[999]);
fulladd full2_439 (sum_2[295], carry_2[295], sum_1[423], carry_1[422], C[1000]);
fulladd full2_440 (sum_2[296], carry_2[296], sum_1[424], carry_1[423], C[1001]);
fulladd full2_441 (sum_2[297], carry_2[297], sum_1[425], carry_1[424], C[1002]);
fulladd full2_442 (sum_2[298], carry_2[298], sum_1[426], carry_1[425], C[1003]);
fulladd full2_443 (sum_2[299], carry_2[299], sum_1[427], carry_1[426], C[1004]);
fulladd full2_444 (sum_2[300], carry_2[300], sum_1[428], carry_1[427], C[1005]);
fulladd full2_445 (sum_2[301], carry_2[301], sum_1[429], carry_1[428], C[1006]);
fulladd full2_446 (sum_2[302], carry_2[302], sum_1[430], carry_1[429], C[1007]);
fulladd full2_447 (sum_2[303], carry_2[303], sum_1[431], carry_1[430], C[1008]);
fulladd full2_448 (sum_2[304], carry_2[304], sum_1[432], carry_1[431], C[1009]);
fulladd full2_449 (sum_2[305], carry_2[305], sum_1[433], carry_1[432], C[1010]);
fulladd full2_450 (sum_2[306], carry_2[306], sum_1[434], carry_1[433], C[1011]);
fulladd full2_451 (sum_2[307], carry_2[307], sum_1[435], carry_1[434], C[1012]);
fulladd full2_452 (sum_2[308], carry_2[308], sum_1[436], carry_1[435], C[1013]);
fulladd full2_453 (sum_2[309], carry_2[309], sum_1[437], carry_1[436], C[1014]);
fulladd full2_454 (sum_2[310], carry_2[310], sum_1[438], carry_1[437], C[1015]);
fulladd full2_455 (sum_2[311], carry_2[311], sum_1[439], carry_1[438], C[1016]);
fulladd full2_456 (sum_2[312], carry_2[312], sum_1[440], carry_1[439], C[1017]);
fulladd full2_457 (sum_2[313], carry_2[313], sum_1[441], carry_1[440], C[1018]);
fulladd full2_458 (sum_2[314], carry_2[314], sum_1[442], carry_1[441], C[1019]);
fulladd full2_459 (sum_2[315], carry_2[315], sum_1[443], carry_1[442], C[1020]);
fulladd full2_460 (sum_2[316], carry_2[316], sum_1[444], carry_1[443], C[1021]);
fulladd full2_461 (sum_2[317], carry_2[317], sum_1[445], carry_1[444], C[1022]);
fulladd full2_462 (sum_2[318], carry_2[318], sum_1[446], carry_1[445], C[1023]);
fulladd full2_463 (sum_2[319], carry_2[319], sum_1[447], carry_1[446], C[1023]);

//sum_2/0/1/2
fulladd full3_00 (sum_3[0], carry_3[0], sum_2[0], sum_2[64], sum_2[128]);
fulladd full3_01 (sum_3[1], carry_3[1], sum_2[1], sum_2[65], sum_2[129]);
fulladd full3_02 (sum_3[2], carry_3[2], sum_2[2], sum_2[66], sum_2[130]);
fulladd full3_03 (sum_3[3], carry_3[3], sum_2[3], sum_2[67], sum_2[131]);
fulladd full3_04 (sum_3[4], carry_3[4], sum_2[4], sum_2[68], sum_2[132]);
fulladd full3_05 (sum_3[5], carry_3[5], sum_2[5], sum_2[69], sum_2[133]);
fulladd full3_06 (sum_3[6], carry_3[6], sum_2[6], sum_2[70], sum_2[134]);
fulladd full3_07 (sum_3[7], carry_3[7], sum_2[7], sum_2[71], sum_2[135]);
fulladd full3_08 (sum_3[8], carry_3[8], sum_2[8], sum_2[72], sum_2[136]);
fulladd full3_09 (sum_3[9], carry_3[9], sum_2[9], sum_2[73], sum_2[137]);
fulladd full3_010 (sum_3[10], carry_3[10], sum_2[10], sum_2[74], sum_2[138]);
fulladd full3_011 (sum_3[11], carry_3[11], sum_2[11], sum_2[75], sum_2[139]);
fulladd full3_012 (sum_3[12], carry_3[12], sum_2[12], sum_2[76], sum_2[140]);
fulladd full3_013 (sum_3[13], carry_3[13], sum_2[13], sum_2[77], sum_2[141]);
fulladd full3_014 (sum_3[14], carry_3[14], sum_2[14], sum_2[78], sum_2[142]);
fulladd full3_015 (sum_3[15], carry_3[15], sum_2[15], sum_2[79], sum_2[143]);
fulladd full3_016 (sum_3[16], carry_3[16], sum_2[16], sum_2[80], sum_2[144]);
fulladd full3_017 (sum_3[17], carry_3[17], sum_2[17], sum_2[81], sum_2[145]);
fulladd full3_018 (sum_3[18], carry_3[18], sum_2[18], sum_2[82], sum_2[146]);
fulladd full3_019 (sum_3[19], carry_3[19], sum_2[19], sum_2[83], sum_2[147]);
fulladd full3_020 (sum_3[20], carry_3[20], sum_2[20], sum_2[84], sum_2[148]);
fulladd full3_021 (sum_3[21], carry_3[21], sum_2[21], sum_2[85], sum_2[149]);
fulladd full3_022 (sum_3[22], carry_3[22], sum_2[22], sum_2[86], sum_2[150]);
fulladd full3_023 (sum_3[23], carry_3[23], sum_2[23], sum_2[87], sum_2[151]);
fulladd full3_024 (sum_3[24], carry_3[24], sum_2[24], sum_2[88], sum_2[152]);
fulladd full3_025 (sum_3[25], carry_3[25], sum_2[25], sum_2[89], sum_2[153]);
fulladd full3_026 (sum_3[26], carry_3[26], sum_2[26], sum_2[90], sum_2[154]);
fulladd full3_027 (sum_3[27], carry_3[27], sum_2[27], sum_2[91], sum_2[155]);
fulladd full3_028 (sum_3[28], carry_3[28], sum_2[28], sum_2[92], sum_2[156]);
fulladd full3_029 (sum_3[29], carry_3[29], sum_2[29], sum_2[93], sum_2[157]);
fulladd full3_030 (sum_3[30], carry_3[30], sum_2[30], sum_2[94], sum_2[158]);
fulladd full3_031 (sum_3[31], carry_3[31], sum_2[31], sum_2[95], sum_2[159]);
fulladd full3_032 (sum_3[32], carry_3[32], sum_2[32], sum_2[96], sum_2[160]);
fulladd full3_033 (sum_3[33], carry_3[33], sum_2[33], sum_2[97], sum_2[161]);
fulladd full3_034 (sum_3[34], carry_3[34], sum_2[34], sum_2[98], sum_2[162]);
fulladd full3_035 (sum_3[35], carry_3[35], sum_2[35], sum_2[99], sum_2[163]);
fulladd full3_036 (sum_3[36], carry_3[36], sum_2[36], sum_2[100], sum_2[164]);
fulladd full3_037 (sum_3[37], carry_3[37], sum_2[37], sum_2[101], sum_2[165]);
fulladd full3_038 (sum_3[38], carry_3[38], sum_2[38], sum_2[102], sum_2[166]);
fulladd full3_039 (sum_3[39], carry_3[39], sum_2[39], sum_2[103], sum_2[167]);
fulladd full3_040 (sum_3[40], carry_3[40], sum_2[40], sum_2[104], sum_2[168]);
fulladd full3_041 (sum_3[41], carry_3[41], sum_2[41], sum_2[105], sum_2[169]);
fulladd full3_042 (sum_3[42], carry_3[42], sum_2[42], sum_2[106], sum_2[170]);
fulladd full3_043 (sum_3[43], carry_3[43], sum_2[43], sum_2[107], sum_2[171]);
fulladd full3_044 (sum_3[44], carry_3[44], sum_2[44], sum_2[108], sum_2[172]);
fulladd full3_045 (sum_3[45], carry_3[45], sum_2[45], sum_2[109], sum_2[173]);
fulladd full3_046 (sum_3[46], carry_3[46], sum_2[46], sum_2[110], sum_2[174]);
fulladd full3_047 (sum_3[47], carry_3[47], sum_2[47], sum_2[111], sum_2[175]);
fulladd full3_048 (sum_3[48], carry_3[48], sum_2[48], sum_2[112], sum_2[176]);
fulladd full3_049 (sum_3[49], carry_3[49], sum_2[49], sum_2[113], sum_2[177]);
fulladd full3_050 (sum_3[50], carry_3[50], sum_2[50], sum_2[114], sum_2[178]);
fulladd full3_051 (sum_3[51], carry_3[51], sum_2[51], sum_2[115], sum_2[179]);
fulladd full3_052 (sum_3[52], carry_3[52], sum_2[52], sum_2[116], sum_2[180]);
fulladd full3_053 (sum_3[53], carry_3[53], sum_2[53], sum_2[117], sum_2[181]);
fulladd full3_054 (sum_3[54], carry_3[54], sum_2[54], sum_2[118], sum_2[182]);
fulladd full3_055 (sum_3[55], carry_3[55], sum_2[55], sum_2[119], sum_2[183]);
fulladd full3_056 (sum_3[56], carry_3[56], sum_2[56], sum_2[120], sum_2[184]);
fulladd full3_057 (sum_3[57], carry_3[57], sum_2[57], sum_2[121], sum_2[185]);
fulladd full3_058 (sum_3[58], carry_3[58], sum_2[58], sum_2[122], sum_2[186]);
fulladd full3_059 (sum_3[59], carry_3[59], sum_2[59], sum_2[123], sum_2[187]);
fulladd full3_060 (sum_3[60], carry_3[60], sum_2[60], sum_2[124], sum_2[188]);
fulladd full3_061 (sum_3[61], carry_3[61], sum_2[61], sum_2[125], sum_2[189]);
fulladd full3_062 (sum_3[62], carry_3[62], sum_2[62], sum_2[126], sum_2[190]);
fulladd full3_063 (sum_3[63], carry_3[63], sum_2[63], sum_2[127], sum_2[191]);

//carry_2/0/1/2
fulladd full3_10 (sum_3[64], carry_3[64], 1'b0, 1'b0, 1'b0);
fulladd full3_11 (sum_3[65], carry_3[65], carry_2[0], carry_2[64], carry_2[128]);
fulladd full3_12 (sum_3[66], carry_3[66], carry_2[1], carry_2[65], carry_2[129]);
fulladd full3_13 (sum_3[67], carry_3[67], carry_2[2], carry_2[66], carry_2[130]);
fulladd full3_14 (sum_3[68], carry_3[68], carry_2[3], carry_2[67], carry_2[131]);
fulladd full3_15 (sum_3[69], carry_3[69], carry_2[4], carry_2[68], carry_2[132]);
fulladd full3_16 (sum_3[70], carry_3[70], carry_2[5], carry_2[69], carry_2[133]);
fulladd full3_17 (sum_3[71], carry_3[71], carry_2[6], carry_2[70], carry_2[134]);
fulladd full3_18 (sum_3[72], carry_3[72], carry_2[7], carry_2[71], carry_2[135]);
fulladd full3_19 (sum_3[73], carry_3[73], carry_2[8], carry_2[72], carry_2[136]);
fulladd full3_110 (sum_3[74], carry_3[74], carry_2[9], carry_2[73], carry_2[137]);
fulladd full3_111 (sum_3[75], carry_3[75], carry_2[10], carry_2[74], carry_2[138]);
fulladd full3_112 (sum_3[76], carry_3[76], carry_2[11], carry_2[75], carry_2[139]);
fulladd full3_113 (sum_3[77], carry_3[77], carry_2[12], carry_2[76], carry_2[140]);
fulladd full3_114 (sum_3[78], carry_3[78], carry_2[13], carry_2[77], carry_2[141]);
fulladd full3_115 (sum_3[79], carry_3[79], carry_2[14], carry_2[78], carry_2[142]);
fulladd full3_116 (sum_3[80], carry_3[80], carry_2[15], carry_2[79], carry_2[143]);
fulladd full3_117 (sum_3[81], carry_3[81], carry_2[16], carry_2[80], carry_2[144]);
fulladd full3_118 (sum_3[82], carry_3[82], carry_2[17], carry_2[81], carry_2[145]);
fulladd full3_119 (sum_3[83], carry_3[83], carry_2[18], carry_2[82], carry_2[146]);
fulladd full3_120 (sum_3[84], carry_3[84], carry_2[19], carry_2[83], carry_2[147]);
fulladd full3_121 (sum_3[85], carry_3[85], carry_2[20], carry_2[84], carry_2[148]);
fulladd full3_122 (sum_3[86], carry_3[86], carry_2[21], carry_2[85], carry_2[149]);
fulladd full3_123 (sum_3[87], carry_3[87], carry_2[22], carry_2[86], carry_2[150]);
fulladd full3_124 (sum_3[88], carry_3[88], carry_2[23], carry_2[87], carry_2[151]);
fulladd full3_125 (sum_3[89], carry_3[89], carry_2[24], carry_2[88], carry_2[152]);
fulladd full3_126 (sum_3[90], carry_3[90], carry_2[25], carry_2[89], carry_2[153]);
fulladd full3_127 (sum_3[91], carry_3[91], carry_2[26], carry_2[90], carry_2[154]);
fulladd full3_128 (sum_3[92], carry_3[92], carry_2[27], carry_2[91], carry_2[155]);
fulladd full3_129 (sum_3[93], carry_3[93], carry_2[28], carry_2[92], carry_2[156]);
fulladd full3_130 (sum_3[94], carry_3[94], carry_2[29], carry_2[93], carry_2[157]);
fulladd full3_131 (sum_3[95], carry_3[95], carry_2[30], carry_2[94], carry_2[158]);
fulladd full3_132 (sum_3[96], carry_3[96], carry_2[31], carry_2[95], carry_2[159]);
fulladd full3_133 (sum_3[97], carry_3[97], carry_2[32], carry_2[96], carry_2[160]);
fulladd full3_134 (sum_3[98], carry_3[98], carry_2[33], carry_2[97], carry_2[161]);
fulladd full3_135 (sum_3[99], carry_3[99], carry_2[34], carry_2[98], carry_2[162]);
fulladd full3_136 (sum_3[100], carry_3[100], carry_2[35], carry_2[99], carry_2[163]);
fulladd full3_137 (sum_3[101], carry_3[101], carry_2[36], carry_2[100], carry_2[164]);
fulladd full3_138 (sum_3[102], carry_3[102], carry_2[37], carry_2[101], carry_2[165]);
fulladd full3_139 (sum_3[103], carry_3[103], carry_2[38], carry_2[102], carry_2[166]);
fulladd full3_140 (sum_3[104], carry_3[104], carry_2[39], carry_2[103], carry_2[167]);
fulladd full3_141 (sum_3[105], carry_3[105], carry_2[40], carry_2[104], carry_2[168]);
fulladd full3_142 (sum_3[106], carry_3[106], carry_2[41], carry_2[105], carry_2[169]);
fulladd full3_143 (sum_3[107], carry_3[107], carry_2[42], carry_2[106], carry_2[170]);
fulladd full3_144 (sum_3[108], carry_3[108], carry_2[43], carry_2[107], carry_2[171]);
fulladd full3_145 (sum_3[109], carry_3[109], carry_2[44], carry_2[108], carry_2[172]);
fulladd full3_146 (sum_3[110], carry_3[110], carry_2[45], carry_2[109], carry_2[173]);
fulladd full3_147 (sum_3[111], carry_3[111], carry_2[46], carry_2[110], carry_2[174]);
fulladd full3_148 (sum_3[112], carry_3[112], carry_2[47], carry_2[111], carry_2[175]);
fulladd full3_149 (sum_3[113], carry_3[113], carry_2[48], carry_2[112], carry_2[176]);
fulladd full3_150 (sum_3[114], carry_3[114], carry_2[49], carry_2[113], carry_2[177]);
fulladd full3_151 (sum_3[115], carry_3[115], carry_2[50], carry_2[114], carry_2[178]);
fulladd full3_152 (sum_3[116], carry_3[116], carry_2[51], carry_2[115], carry_2[179]);
fulladd full3_153 (sum_3[117], carry_3[117], carry_2[52], carry_2[116], carry_2[180]);
fulladd full3_154 (sum_3[118], carry_3[118], carry_2[53], carry_2[117], carry_2[181]);
fulladd full3_155 (sum_3[119], carry_3[119], carry_2[54], carry_2[118], carry_2[182]);
fulladd full3_156 (sum_3[120], carry_3[120], carry_2[55], carry_2[119], carry_2[183]);
fulladd full3_157 (sum_3[121], carry_3[121], carry_2[56], carry_2[120], carry_2[184]);
fulladd full3_158 (sum_3[122], carry_3[122], carry_2[57], carry_2[121], carry_2[185]);
fulladd full3_159 (sum_3[123], carry_3[123], carry_2[58], carry_2[122], carry_2[186]);
fulladd full3_160 (sum_3[124], carry_3[124], carry_2[59], carry_2[123], carry_2[187]);
fulladd full3_161 (sum_3[125], carry_3[125], carry_2[60], carry_2[124], carry_2[188]);
fulladd full3_162 (sum_3[126], carry_3[126], carry_2[61], carry_2[125], carry_2[189]);
fulladd full3_163 (sum_3[127], carry_3[127], carry_2[62], carry_2[126], carry_2[190]);

//sum_2/3/4.carry_3/3
fulladd full3_20 (sum_3[128], carry_3[128], sum_2[192], 1'b0, sum_2[256]);
fulladd full3_21 (sum_3[129], carry_3[129], sum_2[193], carry_2[192], sum_2[257]);
fulladd full3_22 (sum_3[130], carry_3[130], sum_2[194], carry_2[193], sum_2[258]);
fulladd full3_23 (sum_3[131], carry_3[131], sum_2[195], carry_2[194], sum_2[259]);
fulladd full3_24 (sum_3[132], carry_3[132], sum_2[196], carry_2[195], sum_2[260]);
fulladd full3_25 (sum_3[133], carry_3[133], sum_2[197], carry_2[196], sum_2[261]);
fulladd full3_26 (sum_3[134], carry_3[134], sum_2[198], carry_2[197], sum_2[262]);
fulladd full3_27 (sum_3[135], carry_3[135], sum_2[199], carry_2[198], sum_2[263]);
fulladd full3_28 (sum_3[136], carry_3[136], sum_2[200], carry_2[199], sum_2[264]);
fulladd full3_29 (sum_3[137], carry_3[137], sum_2[201], carry_2[200], sum_2[265]);
fulladd full3_210 (sum_3[138], carry_3[138], sum_2[202], carry_2[201], sum_2[266]);
fulladd full3_211 (sum_3[139], carry_3[139], sum_2[203], carry_2[202], sum_2[267]);
fulladd full3_212 (sum_3[140], carry_3[140], sum_2[204], carry_2[203], sum_2[268]);
fulladd full3_213 (sum_3[141], carry_3[141], sum_2[205], carry_2[204], sum_2[269]);
fulladd full3_214 (sum_3[142], carry_3[142], sum_2[206], carry_2[205], sum_2[270]);
fulladd full3_215 (sum_3[143], carry_3[143], sum_2[207], carry_2[206], sum_2[271]);
fulladd full3_216 (sum_3[144], carry_3[144], sum_2[208], carry_2[207], sum_2[272]);
fulladd full3_217 (sum_3[145], carry_3[145], sum_2[209], carry_2[208], sum_2[273]);
fulladd full3_218 (sum_3[146], carry_3[146], sum_2[210], carry_2[209], sum_2[274]);
fulladd full3_219 (sum_3[147], carry_3[147], sum_2[211], carry_2[210], sum_2[275]);
fulladd full3_220 (sum_3[148], carry_3[148], sum_2[212], carry_2[211], sum_2[276]);
fulladd full3_221 (sum_3[149], carry_3[149], sum_2[213], carry_2[212], sum_2[277]);
fulladd full3_222 (sum_3[150], carry_3[150], sum_2[214], carry_2[213], sum_2[278]);
fulladd full3_223 (sum_3[151], carry_3[151], sum_2[215], carry_2[214], sum_2[279]);
fulladd full3_224 (sum_3[152], carry_3[152], sum_2[216], carry_2[215], sum_2[280]);
fulladd full3_225 (sum_3[153], carry_3[153], sum_2[217], carry_2[216], sum_2[281]);
fulladd full3_226 (sum_3[154], carry_3[154], sum_2[218], carry_2[217], sum_2[282]);
fulladd full3_227 (sum_3[155], carry_3[155], sum_2[219], carry_2[218], sum_2[283]);
fulladd full3_228 (sum_3[156], carry_3[156], sum_2[220], carry_2[219], sum_2[284]);
fulladd full3_229 (sum_3[157], carry_3[157], sum_2[221], carry_2[220], sum_2[285]);
fulladd full3_230 (sum_3[158], carry_3[158], sum_2[222], carry_2[221], sum_2[286]);
fulladd full3_231 (sum_3[159], carry_3[159], sum_2[223], carry_2[222], sum_2[287]);
fulladd full3_232 (sum_3[160], carry_3[160], sum_2[224], carry_2[223], sum_2[288]);
fulladd full3_233 (sum_3[161], carry_3[161], sum_2[225], carry_2[224], sum_2[289]);
fulladd full3_234 (sum_3[162], carry_3[162], sum_2[226], carry_2[225], sum_2[290]);
fulladd full3_235 (sum_3[163], carry_3[163], sum_2[227], carry_2[226], sum_2[291]);
fulladd full3_236 (sum_3[164], carry_3[164], sum_2[228], carry_2[227], sum_2[292]);
fulladd full3_237 (sum_3[165], carry_3[165], sum_2[229], carry_2[228], sum_2[293]);
fulladd full3_238 (sum_3[166], carry_3[166], sum_2[230], carry_2[229], sum_2[294]);
fulladd full3_239 (sum_3[167], carry_3[167], sum_2[231], carry_2[230], sum_2[295]);
fulladd full3_240 (sum_3[168], carry_3[168], sum_2[232], carry_2[231], sum_2[296]);
fulladd full3_241 (sum_3[169], carry_3[169], sum_2[233], carry_2[232], sum_2[297]);
fulladd full3_242 (sum_3[170], carry_3[170], sum_2[234], carry_2[233], sum_2[298]);
fulladd full3_243 (sum_3[171], carry_3[171], sum_2[235], carry_2[234], sum_2[299]);
fulladd full3_244 (sum_3[172], carry_3[172], sum_2[236], carry_2[235], sum_2[300]);
fulladd full3_245 (sum_3[173], carry_3[173], sum_2[237], carry_2[236], sum_2[301]);
fulladd full3_246 (sum_3[174], carry_3[174], sum_2[238], carry_2[237], sum_2[302]);
fulladd full3_247 (sum_3[175], carry_3[175], sum_2[239], carry_2[238], sum_2[303]);
fulladd full3_248 (sum_3[176], carry_3[176], sum_2[240], carry_2[239], sum_2[304]);
fulladd full3_249 (sum_3[177], carry_3[177], sum_2[241], carry_2[240], sum_2[305]);
fulladd full3_250 (sum_3[178], carry_3[178], sum_2[242], carry_2[241], sum_2[306]);
fulladd full3_251 (sum_3[179], carry_3[179], sum_2[243], carry_2[242], sum_2[307]);
fulladd full3_252 (sum_3[180], carry_3[180], sum_2[244], carry_2[243], sum_2[308]);
fulladd full3_253 (sum_3[181], carry_3[181], sum_2[245], carry_2[244], sum_2[309]);
fulladd full3_254 (sum_3[182], carry_3[182], sum_2[246], carry_2[245], sum_2[310]);
fulladd full3_255 (sum_3[183], carry_3[183], sum_2[247], carry_2[246], sum_2[311]);
fulladd full3_256 (sum_3[184], carry_3[184], sum_2[248], carry_2[247], sum_2[312]);
fulladd full3_257 (sum_3[185], carry_3[185], sum_2[249], carry_2[248], sum_2[313]);
fulladd full3_258 (sum_3[186], carry_3[186], sum_2[250], carry_2[249], sum_2[314]);
fulladd full3_259 (sum_3[187], carry_3[187], sum_2[251], carry_2[250], sum_2[315]);
fulladd full3_260 (sum_3[188], carry_3[188], sum_2[252], carry_2[251], sum_2[316]);
fulladd full3_261 (sum_3[189], carry_3[189], sum_2[253], carry_2[252], sum_2[317]);
fulladd full3_262 (sum_3[190], carry_3[190], sum_2[254], carry_2[253], sum_2[318]);
fulladd full3_263 (sum_3[191], carry_3[191], sum_2[255], carry_2[254], sum_2[319]);

//sum_3/0/1/2
fulladd full4_00 (sum_4[0], carry_4[0], sum_3[0], sum_3[64], sum_3[128]);
fulladd full4_01 (sum_4[1], carry_4[1], sum_3[1], sum_3[65], sum_3[129]);
fulladd full4_02 (sum_4[2], carry_4[2], sum_3[2], sum_3[66], sum_3[130]);
fulladd full4_03 (sum_4[3], carry_4[3], sum_3[3], sum_3[67], sum_3[131]);
fulladd full4_04 (sum_4[4], carry_4[4], sum_3[4], sum_3[68], sum_3[132]);
fulladd full4_05 (sum_4[5], carry_4[5], sum_3[5], sum_3[69], sum_3[133]);
fulladd full4_06 (sum_4[6], carry_4[6], sum_3[6], sum_3[70], sum_3[134]);
fulladd full4_07 (sum_4[7], carry_4[7], sum_3[7], sum_3[71], sum_3[135]);
fulladd full4_08 (sum_4[8], carry_4[8], sum_3[8], sum_3[72], sum_3[136]);
fulladd full4_09 (sum_4[9], carry_4[9], sum_3[9], sum_3[73], sum_3[137]);
fulladd full4_010 (sum_4[10], carry_4[10], sum_3[10], sum_3[74], sum_3[138]);
fulladd full4_011 (sum_4[11], carry_4[11], sum_3[11], sum_3[75], sum_3[139]);
fulladd full4_012 (sum_4[12], carry_4[12], sum_3[12], sum_3[76], sum_3[140]);
fulladd full4_013 (sum_4[13], carry_4[13], sum_3[13], sum_3[77], sum_3[141]);
fulladd full4_014 (sum_4[14], carry_4[14], sum_3[14], sum_3[78], sum_3[142]);
fulladd full4_015 (sum_4[15], carry_4[15], sum_3[15], sum_3[79], sum_3[143]);
fulladd full4_016 (sum_4[16], carry_4[16], sum_3[16], sum_3[80], sum_3[144]);
fulladd full4_017 (sum_4[17], carry_4[17], sum_3[17], sum_3[81], sum_3[145]);
fulladd full4_018 (sum_4[18], carry_4[18], sum_3[18], sum_3[82], sum_3[146]);
fulladd full4_019 (sum_4[19], carry_4[19], sum_3[19], sum_3[83], sum_3[147]);
fulladd full4_020 (sum_4[20], carry_4[20], sum_3[20], sum_3[84], sum_3[148]);
fulladd full4_021 (sum_4[21], carry_4[21], sum_3[21], sum_3[85], sum_3[149]);
fulladd full4_022 (sum_4[22], carry_4[22], sum_3[22], sum_3[86], sum_3[150]);
fulladd full4_023 (sum_4[23], carry_4[23], sum_3[23], sum_3[87], sum_3[151]);
fulladd full4_024 (sum_4[24], carry_4[24], sum_3[24], sum_3[88], sum_3[152]);
fulladd full4_025 (sum_4[25], carry_4[25], sum_3[25], sum_3[89], sum_3[153]);
fulladd full4_026 (sum_4[26], carry_4[26], sum_3[26], sum_3[90], sum_3[154]);
fulladd full4_027 (sum_4[27], carry_4[27], sum_3[27], sum_3[91], sum_3[155]);
fulladd full4_028 (sum_4[28], carry_4[28], sum_3[28], sum_3[92], sum_3[156]);
fulladd full4_029 (sum_4[29], carry_4[29], sum_3[29], sum_3[93], sum_3[157]);
fulladd full4_030 (sum_4[30], carry_4[30], sum_3[30], sum_3[94], sum_3[158]);
fulladd full4_031 (sum_4[31], carry_4[31], sum_3[31], sum_3[95], sum_3[159]);
fulladd full4_032 (sum_4[32], carry_4[32], sum_3[32], sum_3[96], sum_3[160]);
fulladd full4_033 (sum_4[33], carry_4[33], sum_3[33], sum_3[97], sum_3[161]);
fulladd full4_034 (sum_4[34], carry_4[34], sum_3[34], sum_3[98], sum_3[162]);
fulladd full4_035 (sum_4[35], carry_4[35], sum_3[35], sum_3[99], sum_3[163]);
fulladd full4_036 (sum_4[36], carry_4[36], sum_3[36], sum_3[100], sum_3[164]);
fulladd full4_037 (sum_4[37], carry_4[37], sum_3[37], sum_3[101], sum_3[165]);
fulladd full4_038 (sum_4[38], carry_4[38], sum_3[38], sum_3[102], sum_3[166]);
fulladd full4_039 (sum_4[39], carry_4[39], sum_3[39], sum_3[103], sum_3[167]);
fulladd full4_040 (sum_4[40], carry_4[40], sum_3[40], sum_3[104], sum_3[168]);
fulladd full4_041 (sum_4[41], carry_4[41], sum_3[41], sum_3[105], sum_3[169]);
fulladd full4_042 (sum_4[42], carry_4[42], sum_3[42], sum_3[106], sum_3[170]);
fulladd full4_043 (sum_4[43], carry_4[43], sum_3[43], sum_3[107], sum_3[171]);
fulladd full4_044 (sum_4[44], carry_4[44], sum_3[44], sum_3[108], sum_3[172]);
fulladd full4_045 (sum_4[45], carry_4[45], sum_3[45], sum_3[109], sum_3[173]);
fulladd full4_046 (sum_4[46], carry_4[46], sum_3[46], sum_3[110], sum_3[174]);
fulladd full4_047 (sum_4[47], carry_4[47], sum_3[47], sum_3[111], sum_3[175]);
fulladd full4_048 (sum_4[48], carry_4[48], sum_3[48], sum_3[112], sum_3[176]);
fulladd full4_049 (sum_4[49], carry_4[49], sum_3[49], sum_3[113], sum_3[177]);
fulladd full4_050 (sum_4[50], carry_4[50], sum_3[50], sum_3[114], sum_3[178]);
fulladd full4_051 (sum_4[51], carry_4[51], sum_3[51], sum_3[115], sum_3[179]);
fulladd full4_052 (sum_4[52], carry_4[52], sum_3[52], sum_3[116], sum_3[180]);
fulladd full4_053 (sum_4[53], carry_4[53], sum_3[53], sum_3[117], sum_3[181]);
fulladd full4_054 (sum_4[54], carry_4[54], sum_3[54], sum_3[118], sum_3[182]);
fulladd full4_055 (sum_4[55], carry_4[55], sum_3[55], sum_3[119], sum_3[183]);
fulladd full4_056 (sum_4[56], carry_4[56], sum_3[56], sum_3[120], sum_3[184]);
fulladd full4_057 (sum_4[57], carry_4[57], sum_3[57], sum_3[121], sum_3[185]);
fulladd full4_058 (sum_4[58], carry_4[58], sum_3[58], sum_3[122], sum_3[186]);
fulladd full4_059 (sum_4[59], carry_4[59], sum_3[59], sum_3[123], sum_3[187]);
fulladd full4_060 (sum_4[60], carry_4[60], sum_3[60], sum_3[124], sum_3[188]);
fulladd full4_061 (sum_4[61], carry_4[61], sum_3[61], sum_3[125], sum_3[189]);
fulladd full4_062 (sum_4[62], carry_4[62], sum_3[62], sum_3[126], sum_3[190]);
fulladd full4_063 (sum_4[63], carry_4[63], sum_3[63], sum_3[127], sum_3[191]);

//carry_3/0/1/2
fulladd full4_10 (sum_4[64], carry_4[64], 1'b0, 1'b0, 1'b0);
fulladd full4_11 (sum_4[65], carry_4[65], carry_3[0], carry_3[64], carry_3[128]);
fulladd full4_12 (sum_4[66], carry_4[66], carry_3[1], carry_3[65], carry_3[129]);
fulladd full4_13 (sum_4[67], carry_4[67], carry_3[2], carry_3[66], carry_3[130]);
fulladd full4_14 (sum_4[68], carry_4[68], carry_3[3], carry_3[67], carry_3[131]);
fulladd full4_15 (sum_4[69], carry_4[69], carry_3[4], carry_3[68], carry_3[132]);
fulladd full4_16 (sum_4[70], carry_4[70], carry_3[5], carry_3[69], carry_3[133]);
fulladd full4_17 (sum_4[71], carry_4[71], carry_3[6], carry_3[70], carry_3[134]);
fulladd full4_18 (sum_4[72], carry_4[72], carry_3[7], carry_3[71], carry_3[135]);
fulladd full4_19 (sum_4[73], carry_4[73], carry_3[8], carry_3[72], carry_3[136]);
fulladd full4_110 (sum_4[74], carry_4[74], carry_3[9], carry_3[73], carry_3[137]);
fulladd full4_111 (sum_4[75], carry_4[75], carry_3[10], carry_3[74], carry_3[138]);
fulladd full4_112 (sum_4[76], carry_4[76], carry_3[11], carry_3[75], carry_3[139]);
fulladd full4_113 (sum_4[77], carry_4[77], carry_3[12], carry_3[76], carry_3[140]);
fulladd full4_114 (sum_4[78], carry_4[78], carry_3[13], carry_3[77], carry_3[141]);
fulladd full4_115 (sum_4[79], carry_4[79], carry_3[14], carry_3[78], carry_3[142]);
fulladd full4_116 (sum_4[80], carry_4[80], carry_3[15], carry_3[79], carry_3[143]);
fulladd full4_117 (sum_4[81], carry_4[81], carry_3[16], carry_3[80], carry_3[144]);
fulladd full4_118 (sum_4[82], carry_4[82], carry_3[17], carry_3[81], carry_3[145]);
fulladd full4_119 (sum_4[83], carry_4[83], carry_3[18], carry_3[82], carry_3[146]);
fulladd full4_120 (sum_4[84], carry_4[84], carry_3[19], carry_3[83], carry_3[147]);
fulladd full4_121 (sum_4[85], carry_4[85], carry_3[20], carry_3[84], carry_3[148]);
fulladd full4_122 (sum_4[86], carry_4[86], carry_3[21], carry_3[85], carry_3[149]);
fulladd full4_123 (sum_4[87], carry_4[87], carry_3[22], carry_3[86], carry_3[150]);
fulladd full4_124 (sum_4[88], carry_4[88], carry_3[23], carry_3[87], carry_3[151]);
fulladd full4_125 (sum_4[89], carry_4[89], carry_3[24], carry_3[88], carry_3[152]);
fulladd full4_126 (sum_4[90], carry_4[90], carry_3[25], carry_3[89], carry_3[153]);
fulladd full4_127 (sum_4[91], carry_4[91], carry_3[26], carry_3[90], carry_3[154]);
fulladd full4_128 (sum_4[92], carry_4[92], carry_3[27], carry_3[91], carry_3[155]);
fulladd full4_129 (sum_4[93], carry_4[93], carry_3[28], carry_3[92], carry_3[156]);
fulladd full4_130 (sum_4[94], carry_4[94], carry_3[29], carry_3[93], carry_3[157]);
fulladd full4_131 (sum_4[95], carry_4[95], carry_3[30], carry_3[94], carry_3[158]);
fulladd full4_132 (sum_4[96], carry_4[96], carry_3[31], carry_3[95], carry_3[159]);
fulladd full4_133 (sum_4[97], carry_4[97], carry_3[32], carry_3[96], carry_3[160]);
fulladd full4_134 (sum_4[98], carry_4[98], carry_3[33], carry_3[97], carry_3[161]);
fulladd full4_135 (sum_4[99], carry_4[99], carry_3[34], carry_3[98], carry_3[162]);
fulladd full4_136 (sum_4[100], carry_4[100], carry_3[35], carry_3[99], carry_3[163]);
fulladd full4_137 (sum_4[101], carry_4[101], carry_3[36], carry_3[100], carry_3[164]);
fulladd full4_138 (sum_4[102], carry_4[102], carry_3[37], carry_3[101], carry_3[165]);
fulladd full4_139 (sum_4[103], carry_4[103], carry_3[38], carry_3[102], carry_3[166]);
fulladd full4_140 (sum_4[104], carry_4[104], carry_3[39], carry_3[103], carry_3[167]);
fulladd full4_141 (sum_4[105], carry_4[105], carry_3[40], carry_3[104], carry_3[168]);
fulladd full4_142 (sum_4[106], carry_4[106], carry_3[41], carry_3[105], carry_3[169]);
fulladd full4_143 (sum_4[107], carry_4[107], carry_3[42], carry_3[106], carry_3[170]);
fulladd full4_144 (sum_4[108], carry_4[108], carry_3[43], carry_3[107], carry_3[171]);
fulladd full4_145 (sum_4[109], carry_4[109], carry_3[44], carry_3[108], carry_3[172]);
fulladd full4_146 (sum_4[110], carry_4[110], carry_3[45], carry_3[109], carry_3[173]);
fulladd full4_147 (sum_4[111], carry_4[111], carry_3[46], carry_3[110], carry_3[174]);
fulladd full4_148 (sum_4[112], carry_4[112], carry_3[47], carry_3[111], carry_3[175]);
fulladd full4_149 (sum_4[113], carry_4[113], carry_3[48], carry_3[112], carry_3[176]);
fulladd full4_150 (sum_4[114], carry_4[114], carry_3[49], carry_3[113], carry_3[177]);
fulladd full4_151 (sum_4[115], carry_4[115], carry_3[50], carry_3[114], carry_3[178]);
fulladd full4_152 (sum_4[116], carry_4[116], carry_3[51], carry_3[115], carry_3[179]);
fulladd full4_153 (sum_4[117], carry_4[117], carry_3[52], carry_3[116], carry_3[180]);
fulladd full4_154 (sum_4[118], carry_4[118], carry_3[53], carry_3[117], carry_3[181]);
fulladd full4_155 (sum_4[119], carry_4[119], carry_3[54], carry_3[118], carry_3[182]);
fulladd full4_156 (sum_4[120], carry_4[120], carry_3[55], carry_3[119], carry_3[183]);
fulladd full4_157 (sum_4[121], carry_4[121], carry_3[56], carry_3[120], carry_3[184]);
fulladd full4_158 (sum_4[122], carry_4[122], carry_3[57], carry_3[121], carry_3[185]);
fulladd full4_159 (sum_4[123], carry_4[123], carry_3[58], carry_3[122], carry_3[186]);
fulladd full4_160 (sum_4[124], carry_4[124], carry_3[59], carry_3[123], carry_3[187]);
fulladd full4_161 (sum_4[125], carry_4[125], carry_3[60], carry_3[124], carry_3[188]);
fulladd full4_162 (sum_4[126], carry_4[126], carry_3[61], carry_3[125], carry_3[189]);
fulladd full4_163 (sum_4[127], carry_4[127], carry_3[62], carry_3[126], carry_3[190]);


//sum_4/0/1.carry_4/0
fulladd full5_00 (sum_5[0], carry_5[0], sum_4[0], 1'b0, sum_4[64]);
fulladd full5_01 (sum_5[1], carry_5[1], sum_4[1], carry_4[0], sum_4[65]);
fulladd full5_02 (sum_5[2], carry_5[2], sum_4[2], carry_4[1], sum_4[66]);
fulladd full5_03 (sum_5[3], carry_5[3], sum_4[3], carry_4[2], sum_4[67]);
fulladd full5_04 (sum_5[4], carry_5[4], sum_4[4], carry_4[3], sum_4[68]);
fulladd full5_05 (sum_5[5], carry_5[5], sum_4[5], carry_4[4], sum_4[69]);
fulladd full5_06 (sum_5[6], carry_5[6], sum_4[6], carry_4[5], sum_4[70]);
fulladd full5_07 (sum_5[7], carry_5[7], sum_4[7], carry_4[6], sum_4[71]);
fulladd full5_08 (sum_5[8], carry_5[8], sum_4[8], carry_4[7], sum_4[72]);
fulladd full5_09 (sum_5[9], carry_5[9], sum_4[9], carry_4[8], sum_4[73]);
fulladd full5_010 (sum_5[10], carry_5[10], sum_4[10], carry_4[9], sum_4[74]);
fulladd full5_011 (sum_5[11], carry_5[11], sum_4[11], carry_4[10], sum_4[75]);
fulladd full5_012 (sum_5[12], carry_5[12], sum_4[12], carry_4[11], sum_4[76]);
fulladd full5_013 (sum_5[13], carry_5[13], sum_4[13], carry_4[12], sum_4[77]);
fulladd full5_014 (sum_5[14], carry_5[14], sum_4[14], carry_4[13], sum_4[78]);
fulladd full5_015 (sum_5[15], carry_5[15], sum_4[15], carry_4[14], sum_4[79]);
fulladd full5_016 (sum_5[16], carry_5[16], sum_4[16], carry_4[15], sum_4[80]);
fulladd full5_017 (sum_5[17], carry_5[17], sum_4[17], carry_4[16], sum_4[81]);
fulladd full5_018 (sum_5[18], carry_5[18], sum_4[18], carry_4[17], sum_4[82]);
fulladd full5_019 (sum_5[19], carry_5[19], sum_4[19], carry_4[18], sum_4[83]);
fulladd full5_020 (sum_5[20], carry_5[20], sum_4[20], carry_4[19], sum_4[84]);
fulladd full5_021 (sum_5[21], carry_5[21], sum_4[21], carry_4[20], sum_4[85]);
fulladd full5_022 (sum_5[22], carry_5[22], sum_4[22], carry_4[21], sum_4[86]);
fulladd full5_023 (sum_5[23], carry_5[23], sum_4[23], carry_4[22], sum_4[87]);
fulladd full5_024 (sum_5[24], carry_5[24], sum_4[24], carry_4[23], sum_4[88]);
fulladd full5_025 (sum_5[25], carry_5[25], sum_4[25], carry_4[24], sum_4[89]);
fulladd full5_026 (sum_5[26], carry_5[26], sum_4[26], carry_4[25], sum_4[90]);
fulladd full5_027 (sum_5[27], carry_5[27], sum_4[27], carry_4[26], sum_4[91]);
fulladd full5_028 (sum_5[28], carry_5[28], sum_4[28], carry_4[27], sum_4[92]);
fulladd full5_029 (sum_5[29], carry_5[29], sum_4[29], carry_4[28], sum_4[93]);
fulladd full5_030 (sum_5[30], carry_5[30], sum_4[30], carry_4[29], sum_4[94]);
fulladd full5_031 (sum_5[31], carry_5[31], sum_4[31], carry_4[30], sum_4[95]);
fulladd full5_032 (sum_5[32], carry_5[32], sum_4[32], carry_4[31], sum_4[96]);
fulladd full5_033 (sum_5[33], carry_5[33], sum_4[33], carry_4[32], sum_4[97]);
fulladd full5_034 (sum_5[34], carry_5[34], sum_4[34], carry_4[33], sum_4[98]);
fulladd full5_035 (sum_5[35], carry_5[35], sum_4[35], carry_4[34], sum_4[99]);
fulladd full5_036 (sum_5[36], carry_5[36], sum_4[36], carry_4[35], sum_4[100]);
fulladd full5_037 (sum_5[37], carry_5[37], sum_4[37], carry_4[36], sum_4[101]);
fulladd full5_038 (sum_5[38], carry_5[38], sum_4[38], carry_4[37], sum_4[102]);
fulladd full5_039 (sum_5[39], carry_5[39], sum_4[39], carry_4[38], sum_4[103]);
fulladd full5_040 (sum_5[40], carry_5[40], sum_4[40], carry_4[39], sum_4[104]);
fulladd full5_041 (sum_5[41], carry_5[41], sum_4[41], carry_4[40], sum_4[105]);
fulladd full5_042 (sum_5[42], carry_5[42], sum_4[42], carry_4[41], sum_4[106]);
fulladd full5_043 (sum_5[43], carry_5[43], sum_4[43], carry_4[42], sum_4[107]);
fulladd full5_044 (sum_5[44], carry_5[44], sum_4[44], carry_4[43], sum_4[108]);
fulladd full5_045 (sum_5[45], carry_5[45], sum_4[45], carry_4[44], sum_4[109]);
fulladd full5_046 (sum_5[46], carry_5[46], sum_4[46], carry_4[45], sum_4[110]);
fulladd full5_047 (sum_5[47], carry_5[47], sum_4[47], carry_4[46], sum_4[111]);
fulladd full5_048 (sum_5[48], carry_5[48], sum_4[48], carry_4[47], sum_4[112]);
fulladd full5_049 (sum_5[49], carry_5[49], sum_4[49], carry_4[48], sum_4[113]);
fulladd full5_050 (sum_5[50], carry_5[50], sum_4[50], carry_4[49], sum_4[114]);
fulladd full5_051 (sum_5[51], carry_5[51], sum_4[51], carry_4[50], sum_4[115]);
fulladd full5_052 (sum_5[52], carry_5[52], sum_4[52], carry_4[51], sum_4[116]);
fulladd full5_053 (sum_5[53], carry_5[53], sum_4[53], carry_4[52], sum_4[117]);
fulladd full5_054 (sum_5[54], carry_5[54], sum_4[54], carry_4[53], sum_4[118]);
fulladd full5_055 (sum_5[55], carry_5[55], sum_4[55], carry_4[54], sum_4[119]);
fulladd full5_056 (sum_5[56], carry_5[56], sum_4[56], carry_4[55], sum_4[120]);
fulladd full5_057 (sum_5[57], carry_5[57], sum_4[57], carry_4[56], sum_4[121]);
fulladd full5_058 (sum_5[58], carry_5[58], sum_4[58], carry_4[57], sum_4[122]);
fulladd full5_059 (sum_5[59], carry_5[59], sum_4[59], carry_4[58], sum_4[123]);
fulladd full5_060 (sum_5[60], carry_5[60], sum_4[60], carry_4[59], sum_4[124]);
fulladd full5_061 (sum_5[61], carry_5[61], sum_4[61], carry_4[60], sum_4[125]);
fulladd full5_062 (sum_5[62], carry_5[62], sum_4[62], carry_4[61], sum_4[126]);
fulladd full5_063 (sum_5[63], carry_5[63], sum_4[63], carry_4[62], sum_4[127]);

//sum_5/carry_5/carry_4
fulladd full6_00 (sum_6[0], carry_6[0], sum_5[0], 1'b0, 1'b0);
fulladd full6_01 (sum_6[1], carry_6[1], sum_5[1], carry_5[0], carry_4[64]);
fulladd full6_02 (sum_6[2], carry_6[2], sum_5[2], carry_5[1], carry_4[65]);
fulladd full6_03 (sum_6[3], carry_6[3], sum_5[3], carry_5[2], carry_4[66]);
fulladd full6_04 (sum_6[4], carry_6[4], sum_5[4], carry_5[3], carry_4[67]);
fulladd full6_05 (sum_6[5], carry_6[5], sum_5[5], carry_5[4], carry_4[68]);
fulladd full6_06 (sum_6[6], carry_6[6], sum_5[6], carry_5[5], carry_4[69]);
fulladd full6_07 (sum_6[7], carry_6[7], sum_5[7], carry_5[6], carry_4[70]);
fulladd full6_08 (sum_6[8], carry_6[8], sum_5[8], carry_5[7], carry_4[71]);
fulladd full6_09 (sum_6[9], carry_6[9], sum_5[9], carry_5[8], carry_4[72]);
fulladd full6_010 (sum_6[10], carry_6[10], sum_5[10], carry_5[9], carry_4[73]);
fulladd full6_011 (sum_6[11], carry_6[11], sum_5[11], carry_5[10], carry_4[74]);
fulladd full6_012 (sum_6[12], carry_6[12], sum_5[12], carry_5[11], carry_4[75]);
fulladd full6_013 (sum_6[13], carry_6[13], sum_5[13], carry_5[12], carry_4[76]);
fulladd full6_014 (sum_6[14], carry_6[14], sum_5[14], carry_5[13], carry_4[77]);
fulladd full6_015 (sum_6[15], carry_6[15], sum_5[15], carry_5[14], carry_4[78]);
fulladd full6_016 (sum_6[16], carry_6[16], sum_5[16], carry_5[15], carry_4[79]);
fulladd full6_017 (sum_6[17], carry_6[17], sum_5[17], carry_5[16], carry_4[80]);
fulladd full6_018 (sum_6[18], carry_6[18], sum_5[18], carry_5[17], carry_4[81]);
fulladd full6_019 (sum_6[19], carry_6[19], sum_5[19], carry_5[18], carry_4[82]);
fulladd full6_020 (sum_6[20], carry_6[20], sum_5[20], carry_5[19], carry_4[83]);
fulladd full6_021 (sum_6[21], carry_6[21], sum_5[21], carry_5[20], carry_4[84]);
fulladd full6_022 (sum_6[22], carry_6[22], sum_5[22], carry_5[21], carry_4[85]);
fulladd full6_023 (sum_6[23], carry_6[23], sum_5[23], carry_5[22], carry_4[86]);
fulladd full6_024 (sum_6[24], carry_6[24], sum_5[24], carry_5[23], carry_4[87]);
fulladd full6_025 (sum_6[25], carry_6[25], sum_5[25], carry_5[24], carry_4[88]);
fulladd full6_026 (sum_6[26], carry_6[26], sum_5[26], carry_5[25], carry_4[89]);
fulladd full6_027 (sum_6[27], carry_6[27], sum_5[27], carry_5[26], carry_4[90]);
fulladd full6_028 (sum_6[28], carry_6[28], sum_5[28], carry_5[27], carry_4[91]);
fulladd full6_029 (sum_6[29], carry_6[29], sum_5[29], carry_5[28], carry_4[92]);
fulladd full6_030 (sum_6[30], carry_6[30], sum_5[30], carry_5[29], carry_4[93]);
fulladd full6_031 (sum_6[31], carry_6[31], sum_5[31], carry_5[30], carry_4[94]);
fulladd full6_032 (sum_6[32], carry_6[32], sum_5[32], carry_5[31], carry_4[95]);
fulladd full6_033 (sum_6[33], carry_6[33], sum_5[33], carry_5[32], carry_4[96]);
fulladd full6_034 (sum_6[34], carry_6[34], sum_5[34], carry_5[33], carry_4[97]);
fulladd full6_035 (sum_6[35], carry_6[35], sum_5[35], carry_5[34], carry_4[98]);
fulladd full6_036 (sum_6[36], carry_6[36], sum_5[36], carry_5[35], carry_4[99]);
fulladd full6_037 (sum_6[37], carry_6[37], sum_5[37], carry_5[36], carry_4[100]);
fulladd full6_038 (sum_6[38], carry_6[38], sum_5[38], carry_5[37], carry_4[101]);
fulladd full6_039 (sum_6[39], carry_6[39], sum_5[39], carry_5[38], carry_4[102]);
fulladd full6_040 (sum_6[40], carry_6[40], sum_5[40], carry_5[39], carry_4[103]);
fulladd full6_041 (sum_6[41], carry_6[41], sum_5[41], carry_5[40], carry_4[104]);
fulladd full6_042 (sum_6[42], carry_6[42], sum_5[42], carry_5[41], carry_4[105]);
fulladd full6_043 (sum_6[43], carry_6[43], sum_5[43], carry_5[42], carry_4[106]);
fulladd full6_044 (sum_6[44], carry_6[44], sum_5[44], carry_5[43], carry_4[107]);
fulladd full6_045 (sum_6[45], carry_6[45], sum_5[45], carry_5[44], carry_4[108]);
fulladd full6_046 (sum_6[46], carry_6[46], sum_5[46], carry_5[45], carry_4[109]);
fulladd full6_047 (sum_6[47], carry_6[47], sum_5[47], carry_5[46], carry_4[110]);
fulladd full6_048 (sum_6[48], carry_6[48], sum_5[48], carry_5[47], carry_4[111]);
fulladd full6_049 (sum_6[49], carry_6[49], sum_5[49], carry_5[48], carry_4[112]);
fulladd full6_050 (sum_6[50], carry_6[50], sum_5[50], carry_5[49], carry_4[113]);
fulladd full6_051 (sum_6[51], carry_6[51], sum_5[51], carry_5[50], carry_4[114]);
fulladd full6_052 (sum_6[52], carry_6[52], sum_5[52], carry_5[51], carry_4[115]);
fulladd full6_053 (sum_6[53], carry_6[53], sum_5[53], carry_5[52], carry_4[116]);
fulladd full6_054 (sum_6[54], carry_6[54], sum_5[54], carry_5[53], carry_4[117]);
fulladd full6_055 (sum_6[55], carry_6[55], sum_5[55], carry_5[54], carry_4[118]);
fulladd full6_056 (sum_6[56], carry_6[56], sum_5[56], carry_5[55], carry_4[119]);
fulladd full6_057 (sum_6[57], carry_6[57], sum_5[57], carry_5[56], carry_4[120]);
fulladd full6_058 (sum_6[58], carry_6[58], sum_5[58], carry_5[57], carry_4[121]);
fulladd full6_059 (sum_6[59], carry_6[59], sum_5[59], carry_5[58], carry_4[122]);
fulladd full6_060 (sum_6[60], carry_6[60], sum_5[60], carry_5[59], carry_4[123]);
fulladd full6_061 (sum_6[61], carry_6[61], sum_5[61], carry_5[60], carry_4[124]);
fulladd full6_062 (sum_6[62], carry_6[62], sum_5[62], carry_5[61], carry_4[125]);
fulladd full6_063 (sum_6[63], carry_6[63], sum_5[63], carry_5[62], carry_4[126]);

//sum_6/carry_6/carry_2
fulladd full7_00 (sum_7[0], carry_7[0], sum_6[0], 1'b0, 1'b0);
fulladd full7_01 (sum_7[1], carry_7[1], sum_6[1], carry_6[0], carry_2[256]);
fulladd full7_02 (sum_7[2], carry_7[2], sum_6[2], carry_6[1], carry_2[257]);
fulladd full7_03 (sum_7[3], carry_7[3], sum_6[3], carry_6[2], carry_2[258]);
fulladd full7_04 (sum_7[4], carry_7[4], sum_6[4], carry_6[3], carry_2[259]);
fulladd full7_05 (sum_7[5], carry_7[5], sum_6[5], carry_6[4], carry_2[260]);
fulladd full7_06 (sum_7[6], carry_7[6], sum_6[6], carry_6[5], carry_2[261]);
fulladd full7_07 (sum_7[7], carry_7[7], sum_6[7], carry_6[6], carry_2[262]);
fulladd full7_08 (sum_7[8], carry_7[8], sum_6[8], carry_6[7], carry_2[263]);
fulladd full7_09 (sum_7[9], carry_7[9], sum_6[9], carry_6[8], carry_2[264]);
fulladd full7_010 (sum_7[10], carry_7[10], sum_6[10], carry_6[9], carry_2[265]);
fulladd full7_011 (sum_7[11], carry_7[11], sum_6[11], carry_6[10], carry_2[266]);
fulladd full7_012 (sum_7[12], carry_7[12], sum_6[12], carry_6[11], carry_2[267]);
fulladd full7_013 (sum_7[13], carry_7[13], sum_6[13], carry_6[12], carry_2[268]);
fulladd full7_014 (sum_7[14], carry_7[14], sum_6[14], carry_6[13], carry_2[269]);
fulladd full7_015 (sum_7[15], carry_7[15], sum_6[15], carry_6[14], carry_2[270]);
fulladd full7_016 (sum_7[16], carry_7[16], sum_6[16], carry_6[15], carry_2[271]);
fulladd full7_017 (sum_7[17], carry_7[17], sum_6[17], carry_6[16], carry_2[272]);
fulladd full7_018 (sum_7[18], carry_7[18], sum_6[18], carry_6[17], carry_2[273]);
fulladd full7_019 (sum_7[19], carry_7[19], sum_6[19], carry_6[18], carry_2[274]);
fulladd full7_020 (sum_7[20], carry_7[20], sum_6[20], carry_6[19], carry_2[275]);
fulladd full7_021 (sum_7[21], carry_7[21], sum_6[21], carry_6[20], carry_2[276]);
fulladd full7_022 (sum_7[22], carry_7[22], sum_6[22], carry_6[21], carry_2[277]);
fulladd full7_023 (sum_7[23], carry_7[23], sum_6[23], carry_6[22], carry_2[278]);
fulladd full7_024 (sum_7[24], carry_7[24], sum_6[24], carry_6[23], carry_2[279]);
fulladd full7_025 (sum_7[25], carry_7[25], sum_6[25], carry_6[24], carry_2[280]);
fulladd full7_026 (sum_7[26], carry_7[26], sum_6[26], carry_6[25], carry_2[281]);
fulladd full7_027 (sum_7[27], carry_7[27], sum_6[27], carry_6[26], carry_2[282]);
fulladd full7_028 (sum_7[28], carry_7[28], sum_6[28], carry_6[27], carry_2[283]);
fulladd full7_029 (sum_7[29], carry_7[29], sum_6[29], carry_6[28], carry_2[284]);
fulladd full7_030 (sum_7[30], carry_7[30], sum_6[30], carry_6[29], carry_2[285]);
fulladd full7_031 (sum_7[31], carry_7[31], sum_6[31], carry_6[30], carry_2[286]);
fulladd full7_032 (sum_7[32], carry_7[32], sum_6[32], carry_6[31], carry_2[287]);
fulladd full7_033 (sum_7[33], carry_7[33], sum_6[33], carry_6[32], carry_2[288]);
fulladd full7_034 (sum_7[34], carry_7[34], sum_6[34], carry_6[33], carry_2[289]);
fulladd full7_035 (sum_7[35], carry_7[35], sum_6[35], carry_6[34], carry_2[290]);
fulladd full7_036 (sum_7[36], carry_7[36], sum_6[36], carry_6[35], carry_2[291]);
fulladd full7_037 (sum_7[37], carry_7[37], sum_6[37], carry_6[36], carry_2[292]);
fulladd full7_038 (sum_7[38], carry_7[38], sum_6[38], carry_6[37], carry_2[293]);
fulladd full7_039 (sum_7[39], carry_7[39], sum_6[39], carry_6[38], carry_2[294]);
fulladd full7_040 (sum_7[40], carry_7[40], sum_6[40], carry_6[39], carry_2[295]);
fulladd full7_041 (sum_7[41], carry_7[41], sum_6[41], carry_6[40], carry_2[296]);
fulladd full7_042 (sum_7[42], carry_7[42], sum_6[42], carry_6[41], carry_2[297]);
fulladd full7_043 (sum_7[43], carry_7[43], sum_6[43], carry_6[42], carry_2[298]);
fulladd full7_044 (sum_7[44], carry_7[44], sum_6[44], carry_6[43], carry_2[299]);
fulladd full7_045 (sum_7[45], carry_7[45], sum_6[45], carry_6[44], carry_2[300]);
fulladd full7_046 (sum_7[46], carry_7[46], sum_6[46], carry_6[45], carry_2[301]);
fulladd full7_047 (sum_7[47], carry_7[47], sum_6[47], carry_6[46], carry_2[302]);
fulladd full7_048 (sum_7[48], carry_7[48], sum_6[48], carry_6[47], carry_2[303]);
fulladd full7_049 (sum_7[49], carry_7[49], sum_6[49], carry_6[48], carry_2[304]);
fulladd full7_050 (sum_7[50], carry_7[50], sum_6[50], carry_6[49], carry_2[305]);
fulladd full7_051 (sum_7[51], carry_7[51], sum_6[51], carry_6[50], carry_2[306]);
fulladd full7_052 (sum_7[52], carry_7[52], sum_6[52], carry_6[51], carry_2[307]);
fulladd full7_053 (sum_7[53], carry_7[53], sum_6[53], carry_6[52], carry_2[308]);
fulladd full7_054 (sum_7[54], carry_7[54], sum_6[54], carry_6[53], carry_2[309]);
fulladd full7_055 (sum_7[55], carry_7[55], sum_6[55], carry_6[54], carry_2[310]);
fulladd full7_056 (sum_7[56], carry_7[56], sum_6[56], carry_6[55], carry_2[311]);
fulladd full7_057 (sum_7[57], carry_7[57], sum_6[57], carry_6[56], carry_2[312]);
fulladd full7_058 (sum_7[58], carry_7[58], sum_6[58], carry_6[57], carry_2[313]);
fulladd full7_059 (sum_7[59], carry_7[59], sum_6[59], carry_6[58], carry_2[314]);
fulladd full7_060 (sum_7[60], carry_7[60], sum_6[60], carry_6[59], carry_2[315]);
fulladd full7_061 (sum_7[61], carry_7[61], sum_6[61], carry_6[60], carry_2[316]);
fulladd full7_062 (sum_7[62], carry_7[62], sum_6[62], carry_6[61], carry_2[317]);
fulladd full7_063 (sum_7[63], carry_7[63], sum_6[63], carry_6[62], carry_2[318]);


//final
fulladd full8_00 (O[0], carry_8[0], sum_7[0], 1'b0, 1'b0);
fulladd full8_01 (O[1], carry_8[1], sum_7[1], carry_7[0], carry_8[0]);
fulladd full8_02 (O[2], carry_8[2], sum_7[2], carry_7[1], carry_8[1]);
fulladd full8_03 (O[3], carry_8[3], sum_7[3], carry_7[2], carry_8[2]);
fulladd full8_04 (O[4], carry_8[4], sum_7[4], carry_7[3], carry_8[3]);
fulladd full8_05 (O[5], carry_8[5], sum_7[5], carry_7[4], carry_8[4]);
fulladd full8_06 (O[6], carry_8[6], sum_7[6], carry_7[5], carry_8[5]);
fulladd full8_07 (O[7], carry_8[7], sum_7[7], carry_7[6], carry_8[6]);
fulladd full8_08 (O[8], carry_8[8], sum_7[8], carry_7[7], carry_8[7]);
fulladd full8_09 (O[9], carry_8[9], sum_7[9], carry_7[8], carry_8[8]);
fulladd full8_010 (O[10], carry_8[10], sum_7[10], carry_7[9], carry_8[9]);
fulladd full8_011 (O[11], carry_8[11], sum_7[11], carry_7[10], carry_8[10]);
fulladd full8_012 (O[12], carry_8[12], sum_7[12], carry_7[11], carry_8[11]);
fulladd full8_013 (O[13], carry_8[13], sum_7[13], carry_7[12], carry_8[12]);
fulladd full8_014 (O[14], carry_8[14], sum_7[14], carry_7[13], carry_8[13]);
fulladd full8_015 (O[15], carry_8[15], sum_7[15], carry_7[14], carry_8[14]);
fulladd full8_016 (O[16], carry_8[16], sum_7[16], carry_7[15], carry_8[15]);
fulladd full8_017 (O[17], carry_8[17], sum_7[17], carry_7[16], carry_8[16]);
fulladd full8_018 (O[18], carry_8[18], sum_7[18], carry_7[17], carry_8[17]);
fulladd full8_019 (O[19], carry_8[19], sum_7[19], carry_7[18], carry_8[18]);
fulladd full8_020 (O[20], carry_8[20], sum_7[20], carry_7[19], carry_8[19]);
fulladd full8_021 (O[21], carry_8[21], sum_7[21], carry_7[20], carry_8[20]);
fulladd full8_022 (O[22], carry_8[22], sum_7[22], carry_7[21], carry_8[21]);
fulladd full8_023 (O[23], carry_8[23], sum_7[23], carry_7[22], carry_8[22]);
fulladd full8_024 (O[24], carry_8[24], sum_7[24], carry_7[23], carry_8[23]);
fulladd full8_025 (O[25], carry_8[25], sum_7[25], carry_7[24], carry_8[24]);
fulladd full8_026 (O[26], carry_8[26], sum_7[26], carry_7[25], carry_8[25]);
fulladd full8_027 (O[27], carry_8[27], sum_7[27], carry_7[26], carry_8[26]);
fulladd full8_028 (O[28], carry_8[28], sum_7[28], carry_7[27], carry_8[27]);
fulladd full8_029 (O[29], carry_8[29], sum_7[29], carry_7[28], carry_8[28]);
fulladd full8_030 (O[30], carry_8[30], sum_7[30], carry_7[29], carry_8[29]);
fulladd full8_031 (O[31], carry_8[31], sum_7[31], carry_7[30], carry_8[30]);
fulladd full8_032 (O[32], carry_8[32], sum_7[32], carry_7[31], carry_8[31]);
fulladd full8_033 (O[33], carry_8[33], sum_7[33], carry_7[32], carry_8[32]);
fulladd full8_034 (O[34], carry_8[34], sum_7[34], carry_7[33], carry_8[33]);
fulladd full8_035 (O[35], carry_8[35], sum_7[35], carry_7[34], carry_8[34]);
fulladd full8_036 (O[36], carry_8[36], sum_7[36], carry_7[35], carry_8[35]);
fulladd full8_037 (O[37], carry_8[37], sum_7[37], carry_7[36], carry_8[36]);
fulladd full8_038 (O[38], carry_8[38], sum_7[38], carry_7[37], carry_8[37]);
fulladd full8_039 (O[39], carry_8[39], sum_7[39], carry_7[38], carry_8[38]);
fulladd full8_040 (O[40], carry_8[40], sum_7[40], carry_7[39], carry_8[39]);
fulladd full8_041 (O[41], carry_8[41], sum_7[41], carry_7[40], carry_8[40]);
fulladd full8_042 (O[42], carry_8[42], sum_7[42], carry_7[41], carry_8[41]);
fulladd full8_043 (O[43], carry_8[43], sum_7[43], carry_7[42], carry_8[42]);
fulladd full8_044 (O[44], carry_8[44], sum_7[44], carry_7[43], carry_8[43]);
fulladd full8_045 (O[45], carry_8[45], sum_7[45], carry_7[44], carry_8[44]);
fulladd full8_046 (O[46], carry_8[46], sum_7[46], carry_7[45], carry_8[45]);
fulladd full8_047 (O[47], carry_8[47], sum_7[47], carry_7[46], carry_8[46]);
fulladd full8_048 (O[48], carry_8[48], sum_7[48], carry_7[47], carry_8[47]);
fulladd full8_049 (O[49], carry_8[49], sum_7[49], carry_7[48], carry_8[48]);
fulladd full8_050 (O[50], carry_8[50], sum_7[50], carry_7[49], carry_8[49]);
fulladd full8_051 (O[51], carry_8[51], sum_7[51], carry_7[50], carry_8[50]);
fulladd full8_052 (O[52], carry_8[52], sum_7[52], carry_7[51], carry_8[51]);
fulladd full8_053 (O[53], carry_8[53], sum_7[53], carry_7[52], carry_8[52]);
fulladd full8_054 (O[54], carry_8[54], sum_7[54], carry_7[53], carry_8[53]);
fulladd full8_055 (O[55], carry_8[55], sum_7[55], carry_7[54], carry_8[54]);
fulladd full8_056 (O[56], carry_8[56], sum_7[56], carry_7[55], carry_8[55]);
fulladd full8_057 (O[57], carry_8[57], sum_7[57], carry_7[56], carry_8[56]);
fulladd full8_058 (O[58], carry_8[58], sum_7[58], carry_7[57], carry_8[57]);
fulladd full8_059 (O[59], carry_8[59], sum_7[59], carry_7[58], carry_8[58]);
fulladd full8_060 (O[60], carry_8[60], sum_7[60], carry_7[59], carry_8[59]);
fulladd full8_061 (O[61], carry_8[61], sum_7[61], carry_7[60], carry_8[60]);
fulladd full8_062 (O[62], carry_8[62], sum_7[62], carry_7[61], carry_8[61]);
fulladd full8_063 (O[63], carry_8[63], sum_7[63], carry_7[62], carry_8[62]);

endmodule
