module SDivider(q,r,m,v);
output [31:0]q;
output [31:0]r;
input [31:0]m;
input [31:0]v;
// input [63:0]d;

wire [63:0] d;
wire [31:0] zeros;

assign zeros[31:0] = 0;
assign d[31:0] = v[31:0];
assign d[63:32] = zeros[31:0];

wire [31:0] saksham1, saksham2, saksham3, saksham4, saksham5, saksham6, saksham7, saksham8, saksham9, saksham10, saksham11, saksham12, saksham13, saksham14, saksham15, saksham16, saksham17, saksham18, saksham19, saksham20, saksham21, saksham22, saksham23, saksham24, saksham25, saksham26, saksham27, saksham28, saksham29, saksham30, saksham31, saksham32,saksham33;
wire [31:0]w1;
wire a;
wire [31:0]w2;
wire [31:0]w3;
wire [31:0]w4;
wire [63:0]w5;
wire [31:0]w6;
wire [31:0]s1;
wire [31:0]sum1;
wire [31:0]s2;
wire [31:0]sum2;
wire [31:0]s3;
wire [31:0]sum3;
wire [31:0]s4;
wire [31:0]sum4;
wire [31:0]s5;
wire [31:0]sum5;
wire [31:0]s6;
wire [31:0]sum6;
wire [31:0]s7;
wire [31:0]sum7;
wire [31:0]s8;
wire [31:0]sum8;
wire [31:0]s9;
wire [31:0]sum9;
wire [31:0]s10;
wire [31:0]sum10;
wire [31:0]s11;
wire [31:0]sum11;
wire [31:0]s12;
wire [31:0]sum12;
wire [31:0]s13;
wire [31:0]sum13;
wire [31:0]s14;
wire [31:0]sum14;
wire [31:0]s15;
wire [31:0]sum15;
wire [31:0]s16;
wire [31:0]sum16;
wire [31:0]s17;
wire [31:0]sum17;
wire [31:0]s18;
wire [31:0]sum18;
wire [31:0]s19;
wire [31:0]sum19;
wire [31:0]s20;
wire [31:0]sum20;
wire [31:0]s21;
wire [31:0]sum21;
wire [31:0]s22;
wire [31:0]sum22;
wire [31:0]s23;
wire [31:0]sum23;
wire [31:0]s24;
wire [31:0]sum24;
wire [31:0]s25;
wire [31:0]sum25;
wire [31:0]s26;
wire [31:0]sum26;
wire [31:0]s27;
wire [31:0]sum27;
wire [31:0]s28;
wire [31:0]sum28;
wire [31:0]s29;
wire [31:0]sum29;
wire [31:0]s30;
wire [31:0]sum30;
wire [31:0]s31;
wire [31:0]sum31;
wire [31:0]s32;
wire [31:0]sum32;
wire [31:0]s33;
wire [31:0]sum33;
wire [31:0]sum34;
wire s34;
wire [32:0]q1;
wire [31:0]r1;
wire [32:0]w7;
wire [32:0]w8;
wire [31:0]w9;
wire [31:0]w10;
//converting divisor into normalised form//
xor(w1[31],m[31],m[31]);
xor(w1[30],m[31],m[30]);
xor(w1[29],m[31],m[29]);
xor(w1[28],m[31],m[28]);
xor(w1[27],m[31],m[27]);
xor(w1[26],m[31],m[26]);
xor(w1[25],m[31],m[25]);
xor(w1[24],m[31],m[24]);
xor(w1[23],m[31],m[23]);
xor(w1[22],m[31],m[22]);
xor(w1[21],m[31],m[21]);
xor(w1[20],m[31],m[20]);
xor(w1[19],m[31],m[19]);
xor(w1[18],m[31],m[18]);
xor(w1[17],m[31],m[17]);
xor(w1[16],m[31],m[16]);
xor(w1[15],m[31],m[15]);
xor(w1[14],m[31],m[14]);
xor(w1[13],m[31],m[13]);
xor(w1[12],m[31],m[12]);
xor(w1[11],m[31],m[11]);
xor(w1[10],m[31],m[10]);
xor(w1[9],m[31],m[9]);
xor(w1[8],m[31],m[8]);
xor(w1[7],m[31],m[7]);
xor(w1[6],m[31],m[6]);
xor(w1[5],m[31],m[5]);
xor(w1[4],m[31],m[4]);
xor(w1[3],m[31],m[3]);
xor(w1[2],m[31],m[2]);
xor(w1[1],m[31],m[1]);
xor(w1[0],m[31],m[0]);
//not n6[31:0](r,~w1);

halfadd hd1(w2[0],w3[0],w1[0],m[31]);
halfadd hd2(w2[1],w3[1],w1[1],w3[0]);
halfadd hd3(w2[2],w3[2],w1[2],w3[1]);
halfadd hd4(w2[3],w3[3],w1[3],w3[2]);
halfadd hd5(w2[4],w3[4],w1[4],w3[3]);
halfadd hd6(w2[5],w3[5],w1[5],w3[4]);
halfadd hd7(w2[6],w3[6],w1[6],w3[5]);
halfadd hd8(w2[7],w3[7],w1[7],w3[6]);
halfadd hd9(w2[8],w3[8],w1[8],w3[7]);
halfadd hd10(w2[9],w3[9],w1[9],w3[8]);
halfadd hd11(w2[10],w3[10],w1[10],w3[9]);
halfadd hd12(w2[11],w3[11],w1[11],w3[10]);
halfadd hd13(w2[12],w3[12],w1[12],w3[11]);
halfadd hd14(w2[13],w3[13],w1[13],w3[12]);
halfadd hd15(w2[14],w3[14],w1[14],w3[13]);
halfadd hd16(w2[15],w3[15],w1[15],w3[14]);
halfadd hd17(w2[16],w3[16],w1[16],w3[15]);
halfadd hd18(w2[17],w3[17],w1[17],w3[16]);
halfadd hd19(w2[18],w3[18],w1[18],w3[17]);
halfadd hd20(w2[19],w3[19],w1[19],w3[18]);
halfadd hd21(w2[20],w3[20],w1[20],w3[19]);
halfadd hd22(w2[21],w3[21],w1[21],w3[20]);
halfadd hd23(w2[22],w3[22],w1[22],w3[21]);
halfadd hd24(w2[23],w3[23],w1[23],w3[22]);
halfadd hd25(w2[24],w3[24],w1[24],w3[23]);
halfadd hd26(w2[25],w3[25],w1[25],w3[24]);
halfadd hd27(w2[26],w3[26],w1[26],w3[25]);
halfadd hd28(w2[27],w3[27],w1[27],w3[26]);
halfadd hd29(w2[28],w3[28],w1[28],w3[27]);
halfadd hd30(w2[29],w3[29],w1[29],w3[28]);
halfadd hd31(w2[30],w3[30],w1[30],w3[29]);
halfadd hd32(w2[31],w3[31],w1[31],w3[30]);
//not n6[31:0](r,~w2);

//converting dividend into normalised form//
xor(w4[31],d[31],d[31]);
xor(w4[30],d[31],d[30]);
xor(w4[29],d[31],d[29]);
xor(w4[28],d[31],d[28]);
xor(w4[27],d[31],d[27]);
xor(w4[26],d[31],d[26]);
xor(w4[25],d[31],d[25]);
xor(w4[24],d[31],d[24]);
xor(w4[23],d[31],d[23]);
xor(w4[22],d[31],d[22]);
xor(w4[21],d[31],d[21]);
xor(w4[20],d[31],d[20]);
xor(w4[19],d[31],d[19]);
xor(w4[18],d[31],d[18]);
xor(w4[17],d[31],d[17]);
xor(w4[16],d[31],d[16]);
xor(w4[15],d[31],d[15]);
xor(w4[14],d[31],d[14]);
xor(w4[13],d[31],d[13]);
xor(w4[12],d[31],d[12]);
xor(w4[11],d[31],d[11]);
xor(w4[10],d[31],d[10]);
xor(w4[9],d[31],d[9]);
xor(w4[8],d[31],d[8]);
xor(w4[7],d[31],d[7]);
xor(w4[6],d[31],d[6]);
xor(w4[5],d[31],d[5]);
xor(w4[4],d[31],d[4]);
xor(w4[3],d[31],d[3]);
xor(w4[2],d[31],d[2]);
xor(w4[1],d[31],d[1]);
xor(w4[0],d[31],d[0]);
//not n6[31:0](r,~w4);

halfadd h1(w5[0],w6[0],w4[0],d[31]);
halfadd h2(w5[1],w6[1],w4[1],w6[0]);
halfadd h3(w5[2],w6[2],w4[2],w6[1]);
halfadd h4(w5[3],w6[3],w4[3],w6[2]);
halfadd h5(w5[4],w6[4],w4[4],w6[3]);
halfadd h6(w5[5],w6[5],w4[5],w6[4]);
halfadd h7(w5[6],w6[6],w4[6],w6[5]);
halfadd h8(w5[7],w6[7],w4[7],w6[6]);
halfadd h9(w5[8],w6[8],w4[8],w6[7]);
halfadd h10(w5[9],w6[9],w4[9],w6[8]);
halfadd h11(w5[10],w6[10],w4[10],w6[9]);
halfadd h12(w5[11],w6[11],w4[11],w6[10]);
halfadd h13(w5[12],w6[12],w4[12],w6[11]);
halfadd h14(w5[13],w6[13],w4[13],w6[12]);
halfadd h15(w5[14],w6[14],w4[14],w6[13]);
halfadd h16(w5[15],w6[15],w4[15],w6[14]);
halfadd h17(w5[16],w6[16],w4[16],w6[15]);
halfadd h18(w5[17],w6[17],w4[17],w6[16]);
halfadd h19(w5[18],w6[18],w4[18],w6[17]);
halfadd h20(w5[19],w6[19],w4[19],w6[18]);
halfadd h21(w5[20],w6[20],w4[20],w6[19]);
halfadd h22(w5[21],w6[21],w4[21],w6[20]);
halfadd h23(w5[22],w6[22],w4[22],w6[21]);
halfadd h24(w5[23],w6[23],w4[23],w6[22]);
halfadd h25(w5[24],w6[24],w4[24],w6[23]);
halfadd h26(w5[25],w6[25],w4[25],w3[24]);
halfadd h27(w5[26],w6[26],w4[26],w6[25]);
halfadd h28(w5[27],w6[27],w4[27],w6[26]);
halfadd h29(w5[28],w6[28],w4[28],w6[27]);
halfadd h30(w5[29],w6[29],w4[29],w6[28]);
halfadd h31(w5[30],w6[30],w4[30],w6[29]);
halfadd h32(w5[31],w6[31],w4[31],w6[30]);
//not n6[31:0](r,~w5[31:0]);

//determining sign of quotient and remainder by taking msb bits of divisor and dividend//
xor(a,d[31],m[31]);
//division process//
wire ghj1; 
assign ghj1 = 1;
xor(s1[31],w2[31],ghj1);
xor(s1[30],w2[30],ghj1);
xor(s1[29],w2[29],ghj1);
xor(s1[28],w2[28],ghj1);
xor(s1[27],w2[27],ghj1);
xor(s1[26],w2[26],ghj1);
xor(s1[25],w2[25],ghj1);
xor(s1[24],w2[24],ghj1);
xor(s1[23],w2[23],ghj1);
xor(s1[22],w2[22],ghj1);
xor(s1[21],w2[21],ghj1);
xor(s1[20],w2[20],ghj1);
xor(s1[19],w2[19],ghj1);
xor(s1[18],w2[18],ghj1);
xor(s1[17],w2[17],ghj1);
xor(s1[16],w2[16],ghj1);
xor(s1[15],w2[15],ghj1);
xor(s1[14],w2[14],ghj1);
xor(s1[13],w2[13],ghj1);
xor(s1[12],w2[12],ghj1);
xor(s1[11],w2[11],ghj1);
xor(s1[10],w2[10],ghj1);
xor(s1[9],w2[9],ghj1);
xor(s1[8],w2[8],ghj1);
xor(s1[7],w2[7],ghj1);
xor(s1[6],w2[6],ghj1);
xor(s1[5],w2[5],ghj1);
xor(s1[4],w2[4],ghj1);
xor(s1[3],w2[3],ghj1);
xor(s1[2],w2[2],ghj1);
xor(s1[1],w2[1],ghj1);
xor(s1[0],w2[0],ghj1);

wire ghj; 
assign ghj = 1;
wire [31:0] sehaj,rathore;
//assign sehaj = w5[63:32];
not n2[31:0](w5[63:32],~(32'b0));
assign rathore = s1[31:0];
fulladd32bit fa34(sum1,q1[32],w5[63:32],rathore,ghj);
//not n6(r[0],~q1[32]);


xor(s2[31],w2[31],q1[32]);
xor(s2[30],w2[30],q1[32]);
xor(s2[29],w2[29],q1[32]);
xor(s2[28],w2[28],q1[32]);
xor(s2[27],w2[27],q1[32]);
xor(s2[26],w2[26],q1[32]);
xor(s2[25],w2[25],q1[32]);
xor(s2[24],w2[24],q1[32]);
xor(s2[23],w2[23],q1[32]);
xor(s2[22],w2[22],q1[32]);
xor(s2[21],w2[21],q1[32]);
xor(s2[20],w2[20],q1[32]);
xor(s2[19],w2[19],q1[32]);
xor(s2[18],w2[18],q1[32]);
xor(s2[17],w2[17],q1[32]);
xor(s2[16],w2[16],q1[32]);
xor(s2[15],w2[15],q1[32]);
xor(s2[14],w2[14],q1[32]);
xor(s2[13],w2[13],q1[32]);
xor(s2[12],w2[12],q1[32]);
xor(s2[11],w2[11],q1[32]);
xor(s2[10],w2[10],q1[32]);
xor(s2[9],w2[9],q1[32]);
xor(s2[8],w2[8],q1[32]);
xor(s2[7],w2[7],q1[32]);
xor(s2[6],w2[6],q1[32]);
xor(s2[5],w2[5],q1[32]);
xor(s2[4],w2[4],q1[32]);
xor(s2[3],w2[3],q1[32]);
xor(s2[2],w2[2],q1[32]);
xor(s2[1],w2[1],q1[32]);
xor(s2[0],w2[0],q1[32]);


shifter sh1(saksham1,sum1,w5[31]);
fulladd32bit fa33(sum2,q1[31],saksham1,s2,q1[32]);

xor(s3[31],w2[31],q1[31]);
xor(s3[30],w2[30],q1[31]);
xor(s3[29],w2[29],q1[31]);
xor(s3[28],w2[28],q1[31]);
xor(s3[27],w2[27],q1[31]);
xor(s3[26],w2[26],q1[31]);
xor(s3[25],w2[25],q1[31]);
xor(s3[24],w2[24],q1[31]);
xor(s3[23],w2[23],q1[31]);
xor(s3[22],w2[22],q1[31]);
xor(s3[21],w2[21],q1[31]);
xor(s3[20],w2[20],q1[31]);
xor(s3[19],w2[19],q1[31]);
xor(s3[18],w2[18],q1[31]);
xor(s3[17],w2[17],q1[31]);
xor(s3[16],w2[16],q1[31]);
xor(s3[15],w2[15],q1[31]);
xor(s3[14],w2[14],q1[31]);
xor(s3[13],w2[13],q1[31]);
xor(s3[12],w2[12],q1[31]);
xor(s3[11],w2[11],q1[31]);
xor(s3[10],w2[10],q1[31]);
xor(s3[9],w2[9],q1[31]);
xor(s3[8],w2[8],q1[31]);
xor(s3[7],w2[7],q1[31]);
xor(s3[6],w2[6],q1[31]);
xor(s3[5],w2[5],q1[31]);
xor(s3[4],w2[4],q1[31]);
xor(s3[3],w2[3],q1[31]);
xor(s3[2],w2[2],q1[31]);
xor(s3[1],w2[1],q1[31]);
xor(s3[0],w2[0],q1[31]);


shifter sh2(saksham2,sum2,w5[30]);
fulladd32bit fa32(sum3,q1[30],saksham2,s3,q1[31]);

xor(s4[31],w2[31],q1[30]);
xor(s4[30],w2[30],q1[30]);
xor(s4[29],w2[29],q1[30]);
xor(s4[28],w2[28],q1[30]);
xor(s4[27],w2[27],q1[30]);
xor(s4[26],w2[26],q1[30]);
xor(s4[25],w2[25],q1[30]);
xor(s4[24],w2[24],q1[30]);
xor(s4[23],w2[23],q1[30]);
xor(s4[22],w2[22],q1[30]);
xor(s4[21],w2[21],q1[30]);
xor(s4[20],w2[20],q1[30]);
xor(s4[19],w2[19],q1[30]);
xor(s4[18],w2[18],q1[30]);
xor(s4[17],w2[17],q1[30]);
xor(s4[16],w2[16],q1[30]);
xor(s4[15],w2[15],q1[30]);
xor(s4[14],w2[14],q1[30]);
xor(s4[13],w2[13],q1[30]);
xor(s4[12],w2[12],q1[30]);
xor(s4[11],w2[11],q1[30]);
xor(s4[10],w2[10],q1[30]);
xor(s4[9],w2[9],q1[30]);
xor(s4[8],w2[8],q1[30]);
xor(s4[7],w2[7],q1[30]);
xor(s4[6],w2[6],q1[30]);
xor(s4[5],w2[5],q1[30]);
xor(s4[4],w2[4],q1[30]);
xor(s4[3],w2[3],q1[30]);
xor(s4[2],w2[2],q1[30]);
xor(s4[1],w2[1],q1[30]);
xor(s4[0],w2[0],q1[30]);


shifter sh3(saksham3,sum3,w5[29]);
fulladd32bit fa31(sum4,q1[29],saksham3,s4,q1[30]);

xor(s5[31],w2[31],q1[29]);
xor(s5[30],w2[30],q1[29]);
xor(s5[29],w2[29],q1[29]);
xor(s5[28],w2[28],q1[29]);
xor(s5[27],w2[27],q1[29]);
xor(s5[26],w2[26],q1[29]);
xor(s5[25],w2[25],q1[29]);
xor(s5[24],w2[24],q1[29]);
xor(s5[23],w2[23],q1[29]);
xor(s5[22],w2[22],q1[29]);
xor(s5[21],w2[21],q1[29]);
xor(s5[20],w2[20],q1[29]);
xor(s5[19],w2[19],q1[29]);
xor(s5[18],w2[18],q1[29]);
xor(s5[17],w2[17],q1[29]);
xor(s5[16],w2[16],q1[29]);
xor(s5[15],w2[15],q1[29]);
xor(s5[14],w2[14],q1[29]);
xor(s5[13],w2[13],q1[29]);
xor(s5[12],w2[12],q1[29]);
xor(s5[11],w2[11],q1[29]);
xor(s5[10],w2[10],q1[29]);
xor(s5[9],w2[9],q1[29]);
xor(s5[8],w2[8],q1[29]);
xor(s5[7],w2[7],q1[29]);
xor(s5[6],w2[6],q1[29]);
xor(s5[5],w2[5],q1[29]);
xor(s5[4],w2[4],q1[29]);
xor(s5[3],w2[3],q1[29]);
xor(s5[2],w2[2],q1[29]);
xor(s5[1],w2[1],q1[29]);
xor(s5[0],w2[0],q1[29]);


shifter sh4(saksham4,sum4,w5[28]);
fulladd32bit fa30(sum5,q1[28],saksham4,s5,q1[29]);

xor(s6[31],w2[31],q1[28]);
xor(s6[30],w2[30],q1[28]);
xor(s6[29],w2[29],q1[28]);
xor(s6[28],w2[28],q1[28]);
xor(s6[27],w2[27],q1[28]);
xor(s6[26],w2[26],q1[28]);
xor(s6[25],w2[25],q1[28]);
xor(s6[24],w2[24],q1[28]);
xor(s6[23],w2[23],q1[28]);
xor(s6[22],w2[22],q1[28]);
xor(s6[21],w2[21],q1[28]);
xor(s6[20],w2[20],q1[28]);
xor(s6[19],w2[19],q1[28]);
xor(s6[18],w2[18],q1[28]);
xor(s6[17],w2[17],q1[28]);
xor(s6[16],w2[16],q1[28]);
xor(s6[15],w2[15],q1[28]);
xor(s6[14],w2[14],q1[28]);
xor(s6[13],w2[13],q1[28]);
xor(s6[12],w2[12],q1[28]);
xor(s6[11],w2[11],q1[28]);
xor(s6[10],w2[10],q1[28]);
xor(s6[9],w2[9],q1[28]);
xor(s6[8],w2[8],q1[28]);
xor(s6[7],w2[7],q1[28]);
xor(s6[6],w2[6],q1[28]);
xor(s6[5],w2[5],q1[28]);
xor(s6[4],w2[4],q1[28]);
xor(s6[3],w2[3],q1[28]);
xor(s6[2],w2[2],q1[28]);
xor(s6[1],w2[1],q1[28]);
xor(s6[0],w2[0],q1[28]);


shifter sh5(saksham5,sum5,w5[27]);
fulladd32bit fa29(sum6,q1[27],saksham5,s6,q1[28]);

xor(s7[31],w2[31],q1[27]);
xor(s7[30],w2[30],q1[27]);
xor(s7[29],w2[29],q1[27]);
xor(s7[28],w2[28],q1[27]);
xor(s7[27],w2[27],q1[27]);
xor(s7[26],w2[26],q1[27]);
xor(s7[25],w2[25],q1[27]);
xor(s7[24],w2[24],q1[27]);
xor(s7[23],w2[23],q1[27]);
xor(s7[22],w2[22],q1[27]);
xor(s7[21],w2[21],q1[27]);
xor(s7[20],w2[20],q1[27]);
xor(s7[19],w2[19],q1[27]);
xor(s7[18],w2[18],q1[27]);
xor(s7[17],w2[17],q1[27]);
xor(s7[16],w2[16],q1[27]);
xor(s7[15],w2[15],q1[27]);
xor(s7[14],w2[14],q1[27]);
xor(s7[13],w2[13],q1[27]);
xor(s7[12],w2[12],q1[27]);
xor(s7[11],w2[11],q1[27]);
xor(s7[10],w2[10],q1[27]);
xor(s7[9],w2[9],q1[27]);
xor(s7[8],w2[8],q1[27]);
xor(s7[7],w2[7],q1[27]);
xor(s7[6],w2[6],q1[27]);
xor(s7[5],w2[5],q1[27]);
xor(s7[4],w2[4],q1[27]);
xor(s7[3],w2[3],q1[27]);
xor(s7[2],w2[2],q1[27]);
xor(s7[1],w2[1],q1[27]);
xor(s7[0],w2[0],q1[27]);


shifter sh6(saksham6,sum6,w5[26]);
fulladd32bit fa28(sum7,q1[26],saksham6,s7,q1[27]);


xor(s8[31],w2[31],q1[26]);
xor(s8[30],w2[30],q1[26]);
xor(s8[29],w2[29],q1[26]);
xor(s8[28],w2[28],q1[26]);
xor(s8[27],w2[27],q1[26]);
xor(s8[26],w2[26],q1[26]);
xor(s8[25],w2[25],q1[26]);
xor(s8[24],w2[24],q1[26]);
xor(s8[23],w2[23],q1[26]);
xor(s8[22],w2[22],q1[26]);
xor(s8[21],w2[21],q1[26]);
xor(s8[20],w2[20],q1[26]);
xor(s8[19],w2[19],q1[26]);
xor(s8[18],w2[18],q1[26]);
xor(s8[17],w2[17],q1[26]);
xor(s8[16],w2[16],q1[26]);
xor(s8[15],w2[15],q1[26]);
xor(s8[14],w2[14],q1[26]);
xor(s8[13],w2[13],q1[26]);
xor(s8[12],w2[12],q1[26]);
xor(s8[11],w2[11],q1[26]);
xor(s8[10],w2[10],q1[26]);
xor(s8[9],w2[9],q1[26]);
xor(s8[8],w2[8],q1[26]);
xor(s8[7],w2[7],q1[26]);
xor(s8[6],w2[6],q1[26]);
xor(s8[5],w2[5],q1[26]);
xor(s8[4],w2[4],q1[26]);
xor(s8[3],w2[3],q1[26]);
xor(s8[2],w2[2],q1[26]);
xor(s8[1],w2[1],q1[26]);
xor(s8[0],w2[0],q1[26]);

//not n4[31:0](r,~(s8));
shifter sh7(saksham7,sum7,w5[25]);
fulladd32bit fa27(sum8,q1[25],saksham7,s8,q1[26]);
//not n4[31:0](r,~(sum8));


xor(s9[31],w2[31],q1[25]);
xor(s9[30],w2[30],q1[25]);
xor(s9[29],w2[29],q1[25]);
xor(s9[28],w2[28],q1[25]);
xor(s9[27],w2[27],q1[25]);
xor(s9[26],w2[26],q1[25]);
xor(s9[25],w2[25],q1[25]);
xor(s9[24],w2[24],q1[25]);
xor(s9[23],w2[23],q1[25]);
xor(s9[22],w2[22],q1[25]);
xor(s9[21],w2[21],q1[25]);
xor(s9[20],w2[20],q1[25]);
xor(s9[19],w2[19],q1[25]);
xor(s9[18],w2[18],q1[25]);
xor(s9[17],w2[17],q1[25]);
xor(s9[16],w2[16],q1[25]);
xor(s9[15],w2[15],q1[25]);
xor(s9[14],w2[14],q1[25]);
xor(s9[13],w2[13],q1[25]);
xor(s9[12],w2[12],q1[25]);
xor(s9[11],w2[11],q1[25]);
xor(s9[10],w2[10],q1[25]);
xor(s9[9],w2[9],q1[25]);
xor(s9[8],w2[8],q1[25]);
xor(s9[7],w2[7],q1[25]);
xor(s9[6],w2[6],q1[25]);
xor(s9[5],w2[5],q1[25]);
xor(s9[4],w2[4],q1[25]);
xor(s9[3],w2[3],q1[25]);
xor(s9[2],w2[2],q1[25]);
xor(s9[1],w2[1],q1[25]);
xor(s9[0],w2[0],q1[25]);


shifter sh8(saksham8,sum8,w5[24]);
fulladd32bit fa26(sum9,q1[24],saksham8,s9,q1[25]);

xor(s10[31],w2[31],q1[24]);
xor(s10[30],w2[30],q1[24]);
xor(s10[29],w2[29],q1[24]);
xor(s10[28],w2[28],q1[24]);
xor(s10[27],w2[27],q1[24]);
xor(s10[26],w2[26],q1[24]);
xor(s10[25],w2[25],q1[24]);
xor(s10[24],w2[24],q1[24]);
xor(s10[23],w2[23],q1[24]);
xor(s10[22],w2[22],q1[24]);
xor(s10[21],w2[21],q1[24]);
xor(s10[20],w2[20],q1[24]);
xor(s10[19],w2[19],q1[24]);
xor(s10[18],w2[18],q1[24]);
xor(s10[17],w2[17],q1[24]);
xor(s10[16],w2[16],q1[24]);
xor(s10[15],w2[15],q1[24]);
xor(s10[14],w2[14],q1[24]);
xor(s10[13],w2[13],q1[24]);
xor(s10[12],w2[12],q1[24]);
xor(s10[11],w2[11],q1[24]);
xor(s10[10],w2[10],q1[24]);
xor(s10[9],w2[9],q1[24]);
xor(s10[8],w2[8],q1[24]);
xor(s10[7],w2[7],q1[24]);
xor(s10[6],w2[6],q1[24]);
xor(s10[5],w2[5],q1[24]);
xor(s10[4],w2[4],q1[24]);
xor(s10[3],w2[3],q1[24]);
xor(s10[2],w2[2],q1[24]);
xor(s10[1],w2[1],q1[24]);
xor(s10[0],w2[0],q1[24]);


shifter sh9(saksham9,sum9,w5[23]);
fulladd32bit fa25(sum10,q1[23],saksham9,s10,q1[24]);

xor(s11[31],w2[31],q1[23]);
xor(s11[30],w2[30],q1[23]);
xor(s11[29],w2[29],q1[23]);
xor(s11[28],w2[28],q1[23]);
xor(s11[27],w2[27],q1[23]);
xor(s11[26],w2[26],q1[23]);
xor(s11[25],w2[25],q1[23]);
xor(s11[24],w2[24],q1[23]);
xor(s11[23],w2[23],q1[23]);
xor(s11[22],w2[22],q1[23]);
xor(s11[21],w2[21],q1[23]);
xor(s11[20],w2[20],q1[23]);
xor(s11[19],w2[19],q1[23]);
xor(s11[18],w2[18],q1[23]);
xor(s11[17],w2[17],q1[23]);
xor(s11[16],w2[16],q1[23]);
xor(s11[15],w2[15],q1[23]);
xor(s11[14],w2[14],q1[23]);
xor(s11[13],w2[13],q1[23]);
xor(s11[12],w2[12],q1[23]);
xor(s11[11],w2[11],q1[23]);
xor(s11[10],w2[10],q1[23]);
xor(s11[9],w2[9],q1[23]);
xor(s11[8],w2[8],q1[23]);
xor(s11[7],w2[7],q1[23]);
xor(s11[6],w2[6],q1[23]);
xor(s11[5],w2[5],q1[23]);
xor(s11[4],w2[4],q1[23]);
xor(s11[3],w2[3],q1[23]);
xor(s11[2],w2[2],q1[23]);
xor(s11[1],w2[1],q1[23]);
xor(s11[0],w2[0],q1[23]);


shifter sh10(saksham10,sum10,w5[22]);
fulladd32bit fa24(sum11,q1[22],saksham10,s11,q1[23]);

xor(s12[31],w2[31],q1[22]);
xor(s12[30],w2[30],q1[22]);
xor(s12[29],w2[29],q1[22]);
xor(s12[28],w2[28],q1[22]);
xor(s12[27],w2[27],q1[22]);
xor(s12[26],w2[26],q1[22]);
xor(s12[25],w2[25],q1[22]);
xor(s12[24],w2[24],q1[22]);
xor(s12[23],w2[23],q1[22]);
xor(s12[22],w2[22],q1[22]);
xor(s12[21],w2[21],q1[22]);
xor(s12[20],w2[20],q1[22]);
xor(s12[19],w2[19],q1[22]);
xor(s12[18],w2[18],q1[22]);
xor(s12[17],w2[17],q1[22]);
xor(s12[16],w2[16],q1[22]);
xor(s12[15],w2[15],q1[22]);
xor(s12[14],w2[14],q1[22]);
xor(s12[13],w2[13],q1[22]);
xor(s12[12],w2[12],q1[22]);
xor(s12[11],w2[11],q1[22]);
xor(s12[10],w2[10],q1[22]);
xor(s12[9],w2[9],q1[22]);
xor(s12[8],w2[8],q1[22]);
xor(s12[7],w2[7],q1[22]);
xor(s12[6],w2[6],q1[22]);
xor(s12[5],w2[5],q1[22]);
xor(s12[4],w2[4],q1[22]);
xor(s12[3],w2[3],q1[22]);
xor(s12[2],w2[2],q1[22]);
xor(s12[1],w2[1],q1[22]);
xor(s12[0],w2[0],q1[22]);


shifter sh11(saksham11,sum11,w5[21]);
fulladd32bit fa23(sum12,q1[21],saksham11,s12,q1[22]);

xor(s13[31],w2[31],q1[21]);
xor(s13[30],w2[30],q1[21]);
xor(s13[29],w2[29],q1[21]);
xor(s13[28],w2[28],q1[21]);
xor(s13[27],w2[27],q1[21]);
xor(s13[26],w2[26],q1[21]);
xor(s13[25],w2[25],q1[21]);
xor(s13[24],w2[24],q1[21]);
xor(s13[23],w2[23],q1[21]);
xor(s13[22],w2[22],q1[21]);
xor(s13[21],w2[21],q1[21]);
xor(s13[20],w2[20],q1[21]);
xor(s13[19],w2[19],q1[21]);
xor(s13[18],w2[18],q1[21]);
xor(s13[17],w2[17],q1[21]);
xor(s13[16],w2[16],q1[21]);
xor(s13[15],w2[15],q1[21]);
xor(s13[14],w2[14],q1[21]);
xor(s13[13],w2[13],q1[21]);
xor(s13[12],w2[12],q1[21]);
xor(s13[11],w2[11],q1[21]);
xor(s13[10],w2[10],q1[21]);
xor(s13[9],w2[9],q1[21]);
xor(s13[8],w2[8],q1[21]);
xor(s13[7],w2[7],q1[21]);
xor(s13[6],w2[6],q1[21]);
xor(s13[5],w2[5],q1[21]);
xor(s13[4],w2[4],q1[21]);
xor(s13[3],w2[3],q1[21]);
xor(s13[2],w2[2],q1[21]);
xor(s13[1],w2[1],q1[21]);
xor(s13[0],w2[0],q1[21]);


shifter sh12(saksham12,sum12,w5[20]);
fulladd32bit fa22(sum13,q1[20],saksham12,s13,q1[21]);

xor(s14[31],w2[31],q1[20]);
xor(s14[30],w2[30],q1[20]);
xor(s14[29],w2[29],q1[20]);
xor(s14[28],w2[28],q1[20]);
xor(s14[27],w2[27],q1[20]);
xor(s14[26],w2[26],q1[20]);
xor(s14[25],w2[25],q1[20]);
xor(s14[24],w2[24],q1[20]);
xor(s14[23],w2[23],q1[20]);
xor(s14[22],w2[22],q1[20]);
xor(s14[21],w2[21],q1[20]);
xor(s14[20],w2[20],q1[20]);
xor(s14[19],w2[19],q1[20]);
xor(s14[18],w2[18],q1[20]);
xor(s14[17],w2[17],q1[20]);
xor(s14[16],w2[16],q1[20]);
xor(s14[15],w2[15],q1[20]);
xor(s14[14],w2[14],q1[20]);
xor(s14[13],w2[13],q1[20]);
xor(s14[12],w2[12],q1[20]);
xor(s14[11],w2[11],q1[20]);
xor(s14[10],w2[10],q1[20]);
xor(s14[9],w2[9],q1[20]);
xor(s14[8],w2[8],q1[20]);
xor(s14[7],w2[7],q1[20]);
xor(s14[6],w2[6],q1[20]);
xor(s14[5],w2[5],q1[20]);
xor(s14[4],w2[4],q1[20]);
xor(s14[3],w2[3],q1[20]);
xor(s14[2],w2[2],q1[20]);
xor(s14[1],w2[1],q1[20]);
xor(s14[0],w2[0],q1[20]);


shifter sh13(saksham13,sum13,w5[19]);
fulladd32bit fa21(sum14,q1[19],saksham13,s14,q1[20]);

xor(s15[31],w2[31],q1[19]);
xor(s15[30],w2[30],q1[19]);
xor(s15[29],w2[29],q1[19]);
xor(s15[28],w2[28],q1[19]);
xor(s15[27],w2[27],q1[19]);
xor(s15[26],w2[26],q1[19]);
xor(s15[25],w2[25],q1[19]);
xor(s15[24],w2[24],q1[19]);
xor(s15[23],w2[23],q1[19]);
xor(s15[22],w2[22],q1[19]);
xor(s15[21],w2[21],q1[19]);
xor(s15[20],w2[20],q1[19]);
xor(s15[19],w2[19],q1[19]);
xor(s15[18],w2[18],q1[19]);
xor(s15[17],w2[17],q1[19]);
xor(s15[16],w2[16],q1[19]);
xor(s15[15],w2[15],q1[19]);
xor(s15[14],w2[14],q1[19]);
xor(s15[13],w2[13],q1[19]);
xor(s15[12],w2[12],q1[19]);
xor(s15[11],w2[11],q1[19]);
xor(s15[10],w2[10],q1[19]);
xor(s15[9],w2[9],q1[19]);
xor(s15[8],w2[8],q1[19]);
xor(s15[7],w2[7],q1[19]);
xor(s15[6],w2[6],q1[19]);
xor(s15[5],w2[5],q1[19]);
xor(s15[4],w2[4],q1[19]);
xor(s15[3],w2[3],q1[19]);
xor(s15[2],w2[2],q1[19]);
xor(s15[1],w2[1],q1[19]);
xor(s15[0],w2[0],q1[19]);


shifter sh14(saksham14,sum14,w5[18]);
fulladd32bit fa20(sum15,q1[18],saksham14,s15,q1[19]);

xor(s16[31],w2[31],q1[18]);
xor(s16[30],w2[30],q1[18]);
xor(s16[29],w2[29],q1[18]);
xor(s16[28],w2[28],q1[18]);
xor(s16[27],w2[27],q1[18]);
xor(s16[26],w2[26],q1[18]);
xor(s16[25],w2[25],q1[18]);
xor(s16[24],w2[24],q1[18]);
xor(s16[23],w2[23],q1[18]);
xor(s16[22],w2[22],q1[18]);
xor(s16[21],w2[21],q1[18]);
xor(s16[20],w2[20],q1[18]);
xor(s16[19],w2[19],q1[18]);
xor(s16[18],w2[18],q1[18]);
xor(s16[17],w2[17],q1[18]);
xor(s16[16],w2[16],q1[18]);
xor(s16[15],w2[15],q1[18]);
xor(s16[14],w2[14],q1[18]);
xor(s16[13],w2[13],q1[18]);
xor(s16[12],w2[12],q1[18]);
xor(s16[11],w2[11],q1[18]);
xor(s16[10],w2[10],q1[18]);
xor(s16[9],w2[9],q1[18]);
xor(s16[8],w2[8],q1[18]);
xor(s16[7],w2[7],q1[18]);
xor(s16[6],w2[6],q1[18]);
xor(s16[5],w2[5],q1[18]);
xor(s16[4],w2[4],q1[18]);
xor(s16[3],w2[3],q1[18]);
xor(s16[2],w2[2],q1[18]);
xor(s16[1],w2[1],q1[18]);
xor(s16[0],w2[0],q1[18]);


shifter sh15(saksham15,sum15,w5[17]);
fulladd32bit fa19(sum16,q1[17],saksham15,s16,q1[18]);

xor(s17[31],w2[31],q1[17]);
xor(s17[30],w2[30],q1[17]);
xor(s17[29],w2[29],q1[17]);
xor(s17[28],w2[28],q1[17]);
xor(s17[27],w2[27],q1[17]);
xor(s17[26],w2[26],q1[17]);
xor(s17[25],w2[25],q1[17]);
xor(s17[24],w2[24],q1[17]);
xor(s17[23],w2[23],q1[17]);
xor(s17[22],w2[22],q1[17]);
xor(s17[21],w2[21],q1[17]);
xor(s17[20],w2[20],q1[17]);
xor(s17[19],w2[19],q1[17]);
xor(s17[18],w2[18],q1[17]);
xor(s17[17],w2[17],q1[17]);
xor(s17[16],w2[16],q1[17]);
xor(s17[15],w2[15],q1[17]);
xor(s17[14],w2[14],q1[17]);
xor(s17[13],w2[13],q1[17]);
xor(s17[12],w2[12],q1[17]);
xor(s17[11],w2[11],q1[17]);
xor(s17[10],w2[10],q1[17]);
xor(s17[9],w2[9],q1[17]);
xor(s17[8],w2[8],q1[17]);
xor(s17[7],w2[7],q1[17]);
xor(s17[6],w2[6],q1[17]);
xor(s17[5],w2[5],q1[17]);
xor(s17[4],w2[4],q1[17]);
xor(s17[3],w2[3],q1[17]);
xor(s17[2],w2[2],q1[17]);
xor(s17[1],w2[1],q1[17]);
xor(s17[0],w2[0],q1[17]);


shifter sh16(saksham16,sum16,w5[16]);
fulladd32bit fa18(sum17,q1[16],saksham16,s17,q1[17]);

xor(s18[31],w2[31],q1[16]);
xor(s18[30],w2[30],q1[16]);
xor(s18[29],w2[29],q1[16]);
xor(s18[28],w2[28],q1[16]);
xor(s18[27],w2[27],q1[16]);
xor(s18[26],w2[26],q1[16]);
xor(s18[25],w2[25],q1[16]);
xor(s18[24],w2[24],q1[16]);
xor(s18[23],w2[23],q1[16]);
xor(s18[22],w2[22],q1[16]);
xor(s18[21],w2[21],q1[16]);
xor(s18[20],w2[20],q1[16]);
xor(s18[19],w2[19],q1[16]);
xor(s18[18],w2[18],q1[16]);
xor(s18[17],w2[17],q1[16]);
xor(s18[16],w2[16],q1[16]);
xor(s18[15],w2[15],q1[16]);
xor(s18[14],w2[14],q1[16]);
xor(s18[13],w2[13],q1[16]);
xor(s18[12],w2[12],q1[16]);
xor(s18[11],w2[11],q1[16]);
xor(s18[10],w2[10],q1[16]);
xor(s18[9],w2[9],q1[16]);
xor(s18[8],w2[8],q1[16]);
xor(s18[7],w2[7],q1[16]);
xor(s18[6],w2[6],q1[16]);
xor(s18[5],w2[5],q1[16]);
xor(s18[4],w2[4],q1[16]);
xor(s18[3],w2[3],q1[16]);
xor(s18[2],w2[2],q1[16]);
xor(s18[1],w2[1],q1[16]);
xor(s18[0],w2[0],q1[16]);


shifter sh17(saksham17,sum17,w5[15]);
fulladd32bit fa17(sum18,q1[15],saksham17,s18,q1[16]);

xor(s19[31],w2[31],q1[15]);
xor(s19[30],w2[30],q1[15]);
xor(s19[29],w2[29],q1[15]);
xor(s19[28],w2[28],q1[15]);
xor(s19[27],w2[27],q1[15]);
xor(s19[26],w2[26],q1[15]);
xor(s19[25],w2[25],q1[15]);
xor(s19[24],w2[24],q1[15]);
xor(s19[23],w2[23],q1[15]);
xor(s19[22],w2[22],q1[15]);
xor(s19[21],w2[21],q1[15]);
xor(s19[20],w2[20],q1[15]);
xor(s19[19],w2[19],q1[15]);
xor(s19[18],w2[18],q1[15]);
xor(s19[17],w2[17],q1[15]);
xor(s19[16],w2[16],q1[15]);
xor(s19[15],w2[15],q1[15]);
xor(s19[14],w2[14],q1[15]);
xor(s19[13],w2[13],q1[15]);
xor(s19[12],w2[12],q1[15]);
xor(s19[11],w2[11],q1[15]);
xor(s19[10],w2[10],q1[15]);
xor(s19[9],w2[9],q1[15]);
xor(s19[8],w2[8],q1[15]);
xor(s19[7],w2[7],q1[15]);
xor(s19[6],w2[6],q1[15]);
xor(s19[5],w2[5],q1[15]);
xor(s19[4],w2[4],q1[15]);
xor(s19[3],w2[3],q1[15]);
xor(s19[2],w2[2],q1[15]);
xor(s19[1],w2[1],q1[15]);
xor(s19[0],w2[0],q1[15]);


shifter sh18(saksham18,sum18,w5[14]);
fulladd32bit fa16(sum19,q1[14],saksham18,s19,q1[15]);

xor(s20[31],w2[31],q1[14]);
xor(s20[30],w2[30],q1[14]);
xor(s20[29],w2[29],q1[14]);
xor(s20[28],w2[28],q1[14]);
xor(s20[27],w2[27],q1[14]);
xor(s20[26],w2[26],q1[14]);
xor(s20[25],w2[25],q1[14]);
xor(s20[24],w2[24],q1[14]);
xor(s20[23],w2[23],q1[14]);
xor(s20[22],w2[22],q1[14]);
xor(s20[21],w2[21],q1[14]);
xor(s20[20],w2[20],q1[14]);
xor(s20[19],w2[19],q1[14]);
xor(s20[18],w2[18],q1[14]);
xor(s20[17],w2[17],q1[14]);
xor(s20[16],w2[16],q1[14]);
xor(s20[15],w2[15],q1[14]);
xor(s20[14],w2[14],q1[14]);
xor(s20[13],w2[13],q1[14]);
xor(s20[12],w2[12],q1[14]);
xor(s20[11],w2[11],q1[14]);
xor(s20[10],w2[10],q1[14]);
xor(s20[9],w2[9],q1[14]);
xor(s20[8],w2[8],q1[14]);
xor(s20[7],w2[7],q1[14]);
xor(s20[6],w2[6],q1[14]);
xor(s20[5],w2[5],q1[14]);
xor(s20[4],w2[4],q1[14]);
xor(s20[3],w2[3],q1[14]);
xor(s20[2],w2[2],q1[14]);
xor(s20[1],w2[1],q1[14]);
xor(s20[0],w2[0],q1[14]);


shifter sh19(saksham19,sum19,w5[13]);
fulladd32bit fa15(sum20,q1[13],saksham19,s20,q1[14]);

xor(s21[31],w2[31],q1[13]);
xor(s21[30],w2[30],q1[13]);
xor(s21[29],w2[29],q1[13]);
xor(s21[28],w2[28],q1[13]);
xor(s21[27],w2[27],q1[13]);
xor(s21[26],w2[26],q1[13]);
xor(s21[25],w2[25],q1[13]);
xor(s21[24],w2[24],q1[13]);
xor(s21[23],w2[23],q1[13]);
xor(s21[22],w2[22],q1[13]);
xor(s21[21],w2[21],q1[13]);
xor(s21[20],w2[20],q1[13]);
xor(s21[19],w2[19],q1[13]);
xor(s21[18],w2[18],q1[13]);
xor(s21[17],w2[17],q1[13]);
xor(s21[16],w2[16],q1[13]);
xor(s21[15],w2[15],q1[13]);
xor(s21[14],w2[14],q1[13]);
xor(s21[13],w2[13],q1[13]);
xor(s21[12],w2[12],q1[13]);
xor(s21[11],w2[11],q1[13]);
xor(s21[10],w2[10],q1[13]);
xor(s21[9],w2[9],q1[13]);
xor(s21[8],w2[8],q1[13]);
xor(s21[7],w2[7],q1[13]);
xor(s21[6],w2[6],q1[13]);
xor(s21[5],w2[5],q1[13]);
xor(s21[4],w2[4],q1[13]);
xor(s21[3],w2[3],q1[13]);
xor(s21[2],w2[2],q1[13]);
xor(s21[1],w2[1],q1[13]);
xor(s21[0],w2[0],q1[13]);


shifter sh20(saksham20,sum20,w5[12]);
fulladd32bit fa14(sum21,q1[12],saksham20,s21,q1[13]);

xor(s22[31],w2[31],q1[12]);
xor(s22[30],w2[30],q1[12]);
xor(s22[29],w2[29],q1[12]);
xor(s22[28],w2[28],q1[12]);
xor(s22[27],w2[27],q1[12]);
xor(s22[26],w2[26],q1[12]);
xor(s22[25],w2[25],q1[12]);
xor(s22[24],w2[24],q1[12]);
xor(s22[23],w2[23],q1[12]);
xor(s22[22],w2[22],q1[12]);
xor(s22[21],w2[21],q1[12]);
xor(s22[20],w2[20],q1[12]);
xor(s22[19],w2[19],q1[12]);
xor(s22[18],w2[18],q1[12]);
xor(s22[17],w2[17],q1[12]);
xor(s22[16],w2[16],q1[12]);
xor(s22[15],w2[15],q1[12]);
xor(s22[14],w2[14],q1[12]);
xor(s22[13],w2[13],q1[12]);
xor(s22[12],w2[12],q1[12]);
xor(s22[11],w2[11],q1[12]);
xor(s22[10],w2[10],q1[12]);
xor(s22[9],w2[9],q1[12]);
xor(s22[8],w2[8],q1[12]);
xor(s22[7],w2[7],q1[12]);
xor(s22[6],w2[6],q1[12]);
xor(s22[5],w2[5],q1[12]);
xor(s22[4],w2[4],q1[12]);
xor(s22[3],w2[3],q1[12]);
xor(s22[2],w2[2],q1[12]);
xor(s22[1],w2[1],q1[12]);
xor(s22[0],w2[0],q1[12]);


shifter sh21(saksham21,sum21,w5[11]);
fulladd32bit fa13(sum22,q1[11],saksham21,s22,q1[12]);

xor(s23[31],w2[31],q1[11]);
xor(s23[30],w2[30],q1[11]);
xor(s23[29],w2[29],q1[11]);
xor(s23[28],w2[28],q1[11]);
xor(s23[27],w2[27],q1[11]);
xor(s23[26],w2[26],q1[11]);
xor(s23[25],w2[25],q1[11]);
xor(s23[24],w2[24],q1[11]);
xor(s23[23],w2[23],q1[11]);
xor(s23[22],w2[22],q1[11]);
xor(s23[21],w2[21],q1[11]);
xor(s23[20],w2[20],q1[11]);
xor(s23[19],w2[19],q1[11]);
xor(s23[18],w2[18],q1[11]);
xor(s23[17],w2[17],q1[11]);
xor(s23[16],w2[16],q1[11]);
xor(s23[15],w2[15],q1[11]);
xor(s23[14],w2[14],q1[11]);
xor(s23[13],w2[13],q1[11]);
xor(s23[12],w2[12],q1[11]);
xor(s23[11],w2[11],q1[11]);
xor(s23[10],w2[10],q1[11]);
xor(s23[9],w2[9],q1[11]);
xor(s23[8],w2[8],q1[11]);
xor(s23[7],w2[7],q1[11]);
xor(s23[6],w2[6],q1[11]);
xor(s23[5],w2[5],q1[11]);
xor(s23[4],w2[4],q1[11]);
xor(s23[3],w2[3],q1[11]);
xor(s23[2],w2[2],q1[11]);
xor(s23[1],w2[1],q1[11]);
xor(s23[0],w2[0],q1[11]);


shifter sh22(saksham22,sum22,w5[10]);
fulladd32bit fa12(sum23,q1[10],saksham22,s23,q1[11]);

xor(s24[31],w2[31],q1[10]);
xor(s24[30],w2[30],q1[10]);
xor(s24[29],w2[29],q1[10]);
xor(s24[28],w2[28],q1[10]);
xor(s24[27],w2[27],q1[10]);
xor(s24[26],w2[26],q1[10]);
xor(s24[25],w2[25],q1[10]);
xor(s24[24],w2[24],q1[10]);
xor(s24[23],w2[23],q1[10]);
xor(s24[22],w2[22],q1[10]);
xor(s24[21],w2[21],q1[10]);
xor(s24[20],w2[20],q1[10]);
xor(s24[19],w2[19],q1[10]);
xor(s24[18],w2[18],q1[10]);
xor(s24[17],w2[17],q1[10]);
xor(s24[16],w2[16],q1[10]);
xor(s24[15],w2[15],q1[10]);
xor(s24[14],w2[14],q1[10]);
xor(s24[13],w2[13],q1[10]);
xor(s24[12],w2[12],q1[10]);
xor(s24[11],w2[11],q1[10]);
xor(s24[10],w2[10],q1[10]);
xor(s24[9],w2[9],q1[10]);
xor(s24[8],w2[8],q1[10]);
xor(s24[7],w2[7],q1[10]);
xor(s24[6],w2[6],q1[10]);
xor(s24[5],w2[5],q1[10]);
xor(s24[4],w2[4],q1[10]);
xor(s24[3],w2[3],q1[10]);
xor(s24[2],w2[2],q1[10]);
xor(s24[1],w2[1],q1[10]);
xor(s24[0],w2[0],q1[10]);


shifter sh23(saksham23,sum23,w5[9]);
fulladd32bit fa11(sum24,q1[9],saksham23,s24,q1[10]);

xor(s25[31],w2[31],q1[9]);
xor(s25[30],w2[30],q1[9]);
xor(s25[29],w2[29],q1[9]);
xor(s25[28],w2[28],q1[9]);
xor(s25[27],w2[27],q1[9]);
xor(s25[26],w2[26],q1[9]);
xor(s25[25],w2[25],q1[9]);
xor(s25[24],w2[24],q1[9]);
xor(s25[23],w2[23],q1[9]);
xor(s25[22],w2[22],q1[9]);
xor(s25[21],w2[21],q1[9]);
xor(s25[20],w2[20],q1[9]);
xor(s25[19],w2[19],q1[9]);
xor(s25[18],w2[18],q1[9]);
xor(s25[17],w2[17],q1[9]);
xor(s25[16],w2[16],q1[9]);
xor(s25[15],w2[15],q1[9]);
xor(s25[14],w2[14],q1[9]);
xor(s25[13],w2[13],q1[9]);
xor(s25[12],w2[12],q1[9]);
xor(s25[11],w2[11],q1[9]);
xor(s25[10],w2[10],q1[9]);
xor(s25[9],w2[9],q1[9]);
xor(s25[8],w2[8],q1[9]);
xor(s25[7],w2[7],q1[9]);
xor(s25[6],w2[6],q1[9]);
xor(s25[5],w2[5],q1[9]);
xor(s25[4],w2[4],q1[9]);
xor(s25[3],w2[3],q1[9]);
xor(s25[2],w2[2],q1[9]);
xor(s25[1],w2[1],q1[9]);
xor(s25[0],w2[0],q1[9]);


shifter sh24(saksham24,sum24,w5[8]);
fulladd32bit fa10(sum25,q1[8],saksham24,s25,q1[9]);

xor(s26[31],w2[31],q1[8]);
xor(s26[30],w2[30],q1[8]);
xor(s26[29],w2[29],q1[8]);
xor(s26[28],w2[28],q1[8]);
xor(s26[27],w2[27],q1[8]);
xor(s26[26],w2[26],q1[8]);
xor(s26[25],w2[25],q1[8]);
xor(s26[24],w2[24],q1[8]);
xor(s26[23],w2[23],q1[8]);
xor(s26[22],w2[22],q1[8]);
xor(s26[21],w2[21],q1[8]);
xor(s26[20],w2[20],q1[8]);
xor(s26[19],w2[19],q1[8]);
xor(s26[18],w2[18],q1[8]);
xor(s26[17],w2[17],q1[8]);
xor(s26[16],w2[16],q1[8]);
xor(s26[15],w2[15],q1[8]);
xor(s26[14],w2[14],q1[8]);
xor(s26[13],w2[13],q1[8]);
xor(s26[12],w2[12],q1[8]);
xor(s26[11],w2[11],q1[8]);
xor(s26[10],w2[10],q1[8]);
xor(s26[9],w2[9],q1[8]);
xor(s26[8],w2[8],q1[8]);
xor(s26[7],w2[7],q1[8]);
xor(s26[6],w2[6],q1[8]);
xor(s26[5],w2[5],q1[8]);
xor(s26[4],w2[4],q1[8]);
xor(s26[3],w2[3],q1[8]);
xor(s26[2],w2[2],q1[8]);
xor(s26[1],w2[1],q1[8]);
xor(s26[0],w2[0],q1[8]);


shifter sh25(saksham25,sum25,w5[7]);
fulladd32bit fa9(sum26,q1[7],saksham25,s26,q1[8]);

xor(s27[31],w2[31],q1[7]);
xor(s27[30],w2[30],q1[7]);
xor(s27[29],w2[29],q1[7]);
xor(s27[28],w2[28],q1[7]);
xor(s27[27],w2[27],q1[7]);
xor(s27[26],w2[26],q1[7]);
xor(s27[25],w2[25],q1[7]);
xor(s27[24],w2[24],q1[7]);
xor(s27[23],w2[23],q1[7]);
xor(s27[22],w2[22],q1[7]);
xor(s27[21],w2[21],q1[7]);
xor(s27[20],w2[20],q1[7]);
xor(s27[19],w2[19],q1[7]);
xor(s27[18],w2[18],q1[7]);
xor(s27[17],w2[17],q1[7]);
xor(s27[16],w2[16],q1[7]);
xor(s27[15],w2[15],q1[7]);
xor(s27[14],w2[14],q1[7]);
xor(s27[13],w2[13],q1[7]);
xor(s27[12],w2[12],q1[7]);
xor(s27[11],w2[11],q1[7]);
xor(s27[10],w2[10],q1[7]);
xor(s27[9],w2[9],q1[7]);
xor(s27[8],w2[8],q1[7]);
xor(s27[7],w2[7],q1[7]);
xor(s27[6],w2[6],q1[7]);
xor(s27[5],w2[5],q1[7]);
xor(s27[4],w2[4],q1[7]);
xor(s27[3],w2[3],q1[7]);
xor(s27[2],w2[2],q1[7]);
xor(s27[1],w2[1],q1[7]);
xor(s27[0],w2[0],q1[7]);


shifter sh26(saksham26,sum26,w5[6]);
fulladd32bit fa8(sum27,q1[6],saksham26,s27,q1[7]);

xor(s28[31],w2[31],q1[6]);
xor(s28[30],w2[30],q1[6]);
xor(s28[29],w2[29],q1[6]);
xor(s28[28],w2[28],q1[6]);
xor(s28[27],w2[27],q1[6]);
xor(s28[26],w2[26],q1[6]);
xor(s28[25],w2[25],q1[6]);
xor(s28[24],w2[24],q1[6]);
xor(s28[23],w2[23],q1[6]);
xor(s28[22],w2[22],q1[6]);
xor(s28[21],w2[21],q1[6]);
xor(s28[20],w2[20],q1[6]);
xor(s28[19],w2[19],q1[6]);
xor(s28[18],w2[18],q1[6]);
xor(s28[17],w2[17],q1[6]);
xor(s28[16],w2[16],q1[6]);
xor(s28[15],w2[15],q1[6]);
xor(s28[14],w2[14],q1[6]);
xor(s28[13],w2[13],q1[6]);
xor(s28[12],w2[12],q1[6]);
xor(s28[11],w2[11],q1[6]);
xor(s28[10],w2[10],q1[6]);
xor(s28[9],w2[9],q1[6]);
xor(s28[8],w2[8],q1[6]);
xor(s28[7],w2[7],q1[6]);
xor(s28[6],w2[6],q1[6]);
xor(s28[5],w2[5],q1[6]);
xor(s28[4],w2[4],q1[6]);
xor(s28[3],w2[3],q1[6]);
xor(s28[2],w2[2],q1[6]);
xor(s28[1],w2[1],q1[6]);
xor(s28[0],w2[0],q1[6]);


shifter sh27(saksham27,sum27,w5[5]);
fulladd32bit fa7(sum28,q1[5],saksham27,s28,q1[6]);

xor(s29[31],w2[31],q1[5]);
xor(s29[30],w2[30],q1[5]);
xor(s29[29],w2[29],q1[5]);
xor(s29[28],w2[28],q1[5]);
xor(s29[27],w2[27],q1[5]);
xor(s29[26],w2[26],q1[5]);
xor(s29[25],w2[25],q1[5]);
xor(s29[24],w2[24],q1[5]);
xor(s29[23],w2[23],q1[5]);
xor(s29[22],w2[22],q1[5]);
xor(s29[21],w2[21],q1[5]);
xor(s29[20],w2[20],q1[5]);
xor(s29[19],w2[19],q1[5]);
xor(s29[18],w2[18],q1[5]);
xor(s29[17],w2[17],q1[5]);
xor(s29[16],w2[16],q1[5]);
xor(s29[15],w2[15],q1[5]);
xor(s29[14],w2[14],q1[5]);
xor(s29[13],w2[13],q1[5]);
xor(s29[12],w2[12],q1[5]);
xor(s29[11],w2[11],q1[5]);
xor(s29[10],w2[10],q1[5]);
xor(s29[9],w2[9],q1[5]);
xor(s29[8],w2[8],q1[5]);
xor(s29[7],w2[7],q1[5]);
xor(s29[6],w2[6],q1[5]);
xor(s29[5],w2[5],q1[5]);
xor(s29[4],w2[4],q1[5]);
xor(s29[3],w2[3],q1[5]);
xor(s29[2],w2[2],q1[5]);
xor(s29[1],w2[1],q1[5]);
xor(s29[0],w2[0],q1[5]);


shifter sh28(saksham28,sum28,w5[4]);
fulladd32bit fa6(sum29,q1[4],saksham28,s29,q1[5]);

xor(s30[31],w2[31],q1[4]);
xor(s30[30],w2[30],q1[4]);
xor(s30[29],w2[29],q1[4]);
xor(s30[28],w2[28],q1[4]);
xor(s30[27],w2[27],q1[4]);
xor(s30[26],w2[26],q1[4]);
xor(s30[25],w2[25],q1[4]);
xor(s30[24],w2[24],q1[4]);
xor(s30[23],w2[23],q1[4]);
xor(s30[22],w2[22],q1[4]);
xor(s30[21],w2[21],q1[4]);
xor(s30[20],w2[20],q1[4]);
xor(s30[19],w2[19],q1[4]);
xor(s30[18],w2[18],q1[4]);
xor(s30[17],w2[17],q1[4]);
xor(s30[16],w2[16],q1[4]);
xor(s30[15],w2[15],q1[4]);
xor(s30[14],w2[14],q1[4]);
xor(s30[13],w2[13],q1[4]);
xor(s30[12],w2[12],q1[4]);
xor(s30[11],w2[11],q1[4]);
xor(s30[10],w2[10],q1[4]);
xor(s30[9],w2[9],q1[4]);
xor(s30[8],w2[8],q1[4]);
xor(s30[7],w2[7],q1[4]);
xor(s30[6],w2[6],q1[4]);
xor(s30[5],w2[5],q1[4]);
xor(s30[4],w2[4],q1[4]);
xor(s30[3],w2[3],q1[4]);
xor(s30[2],w2[2],q1[4]);
xor(s30[1],w2[1],q1[4]);
xor(s30[0],w2[0],q1[4]);


shifter sh29(saksham29,sum29,w5[3]);
fulladd32bit fa5(sum30,q1[3],saksham29,s30,q1[4]);

xor(s31[31],w2[31],q1[3]);
xor(s31[30],w2[30],q1[3]);
xor(s31[29],w2[29],q1[3]);
xor(s31[28],w2[28],q1[3]);
xor(s31[27],w2[27],q1[3]);
xor(s31[26],w2[26],q1[3]);
xor(s31[25],w2[25],q1[3]);
xor(s31[24],w2[24],q1[3]);
xor(s31[23],w2[23],q1[3]);
xor(s31[22],w2[22],q1[3]);
xor(s31[21],w2[21],q1[3]);
xor(s31[20],w2[20],q1[3]);
xor(s31[19],w2[19],q1[3]);
xor(s31[18],w2[18],q1[3]);
xor(s31[17],w2[17],q1[3]);
xor(s31[16],w2[16],q1[3]);
xor(s31[15],w2[15],q1[3]);
xor(s31[14],w2[14],q1[3]);
xor(s31[13],w2[13],q1[3]);
xor(s31[12],w2[12],q1[3]);
xor(s31[11],w2[11],q1[3]);
xor(s31[10],w2[10],q1[3]);
xor(s31[9],w2[9],q1[3]);
xor(s31[8],w2[8],q1[3]);
xor(s31[7],w2[7],q1[3]);
xor(s31[6],w2[6],q1[3]);
xor(s31[5],w2[5],q1[3]);
xor(s31[4],w2[4],q1[3]);
xor(s31[3],w2[3],q1[3]);
xor(s31[2],w2[2],q1[3]);
xor(s31[1],w2[1],q1[3]);
xor(s31[0],w2[0],q1[3]);


shifter sh30(saksham30,sum30,w5[2]);
fulladd32bit fa4(sum31,q1[2],saksham30,s31,q1[3]);

xor(s32[31],w2[31],q1[2]);
xor(s32[30],w2[30],q1[2]);
xor(s32[29],w2[29],q1[2]);
xor(s32[28],w2[28],q1[2]);
xor(s32[27],w2[27],q1[2]);
xor(s32[26],w2[26],q1[2]);
xor(s32[25],w2[25],q1[2]);
xor(s32[24],w2[24],q1[2]);
xor(s32[23],w2[23],q1[2]);
xor(s32[22],w2[22],q1[2]);
xor(s32[21],w2[21],q1[2]);
xor(s32[20],w2[20],q1[2]);
xor(s32[19],w2[19],q1[2]);
xor(s32[18],w2[18],q1[2]);
xor(s32[17],w2[17],q1[2]);
xor(s32[16],w2[16],q1[2]);
xor(s32[15],w2[15],q1[2]);
xor(s32[14],w2[14],q1[2]);
xor(s32[13],w2[13],q1[2]);
xor(s32[12],w2[12],q1[2]);
xor(s32[11],w2[11],q1[2]);
xor(s32[10],w2[10],q1[2]);
xor(s32[9],w2[9],q1[2]);
xor(s32[8],w2[8],q1[2]);
xor(s32[7],w2[7],q1[2]);
xor(s32[6],w2[6],q1[2]);
xor(s32[5],w2[5],q1[2]);
xor(s32[4],w2[4],q1[2]);
xor(s32[3],w2[3],q1[2]);
xor(s32[2],w2[2],q1[2]);
xor(s32[1],w2[1],q1[2]);
xor(s32[0],w2[0],q1[2]);


shifter sh31(saksham31,sum31,w5[1]);
fulladd32bit fa3(sum32,q1[1], saksham31, s32, q1[2]);

xor(s33[31],w2[31],q1[1]);
xor(s33[30],w2[30],q1[1]);
xor(s33[29],w2[29],q1[1]);
xor(s33[28],w2[28],q1[1]);
xor(s33[27],w2[27],q1[1]);
xor(s33[26],w2[26],q1[1]);
xor(s33[25],w2[25],q1[1]);
xor(s33[24],w2[24],q1[1]);
xor(s33[23],w2[23],q1[1]);
xor(s33[22],w2[22],q1[1]);
xor(s33[21],w2[21],q1[1]);
xor(s33[20],w2[20],q1[1]);
xor(s33[19],w2[19],q1[1]);
xor(s33[18],w2[18],q1[1]);
xor(s33[17],w2[17],q1[1]);
xor(s33[16],w2[16],q1[1]);
xor(s33[15],w2[15],q1[1]);
xor(s33[14],w2[14],q1[1]);
xor(s33[13],w2[13],q1[1]);
xor(s33[12],w2[12],q1[1]);
xor(s33[11],w2[11],q1[1]);
xor(s33[10],w2[10],q1[1]);
xor(s33[9],w2[9],q1[1]);
xor(s33[8],w2[8],q1[1]);
xor(s33[7],w2[7],q1[1]);
xor(s33[6],w2[6],q1[1]);
xor(s33[5],w2[5],q1[1]);
xor(s33[4],w2[4],q1[1]);
xor(s33[3],w2[3],q1[1]);
xor(s33[2],w2[2],q1[1]);
xor(s33[1],w2[1],q1[1]);
xor(s33[0],w2[0],q1[1]);

wire ghj2;
assign ghj2=0;
shifter sh32(saksham32,sum32,w5[0]);
assign saksham33= w2[31:0];
fulladd32bit fa2(sum33,q1[0],saksham32,s33,q1[1]);
fulladd32bit fa1(sum34,s34,sum33,saksham33,ghj2);
mux mx31(r1[31],sum33[31],sum34[31],sum33[31]);
mux mx30(r1[30],sum33[30],sum34[30],sum33[31]);
mux mx29(r1[29],sum33[29],sum34[29],sum33[31]);
mux mx28(r1[28],sum33[28],sum34[28],sum33[31]);
mux mx27(r1[27],sum33[27],sum34[27],sum33[31]);
mux mx26(r1[26],sum33[26],sum34[26],sum33[31]);
mux mx25(r1[25],sum33[25],sum34[25],sum33[31]);
mux mx24(r1[24],sum33[24],sum34[24],sum33[31]);
mux mx23(r1[23],sum33[23],sum34[23],sum33[31]);
mux mx22(r1[22],sum33[22],sum34[22],sum33[31]);
mux mx21(r1[21],sum33[21],sum34[21],sum33[31]);
mux mx20(r1[20],sum33[20],sum34[20],sum33[31]);
mux mx19(r1[19],sum33[19],sum34[19],sum33[31]);
mux mx18(r1[18],sum33[18],sum34[18],sum33[31]);
mux mx17(r1[17],sum33[17],sum34[17],sum33[31]);
mux mx16(r1[16],sum33[16],sum34[16],sum33[31]);
mux mx15(r1[15],sum33[15],sum34[15],sum33[31]);
mux mx14(r1[14],sum33[14],sum34[14],sum33[31]);
mux mx13(r1[13],sum33[13],sum34[13],sum33[31]);
mux mx12(r1[12],sum33[12],sum34[12],sum33[31]);
mux mx11(r1[11],sum33[11],sum34[11],sum33[31]);
mux mx10(r1[10],sum33[10],sum34[10],sum33[31]);
mux mx9(r1[9],sum33[9],sum34[9],sum33[31]);
mux mx8(r1[8],sum33[8],sum34[8],sum33[31]);
mux mx7(r1[7],sum33[7],sum34[7],sum33[31]);
mux mx6(r1[6],sum33[6],sum34[6],sum33[31]);
mux mx5(r1[5],sum33[5],sum34[5],sum33[31]);
mux mx4(r1[4],sum33[4],sum34[4],sum33[31]);
mux mx3(r1[3],sum33[3],sum34[3],sum33[31]);
mux mx2(r1[2],sum33[2],sum34[2],sum33[31]);
mux mx1(r1[1],sum33[1],sum34[1],sum33[31]);
mux mx0(r1[0],sum33[0],sum34[0],sum33[31]);
//not n6[31:0](r,~r1);
//not n6[31:0](r,~q1[31:0]);

//converting normalised form of quotient into output form//

//xor(w7[32],a,q1[32]);
//not n6(r[0],~w7[32]);

xor(w7[31],a,q1[31]);
//not n6(r[0],~w7[31]);
xor(w7[30],a,q1[30]);
xor(w7[29],a,q1[29]);
xor(w7[28],a,q1[28]);
xor(w7[27],a,q1[27]);
xor(w7[26],a,q1[26]);
xor(w7[25],a,q1[25]);
xor(w7[24],a,q1[24]);
xor(w7[23],a,q1[23]);
xor(w7[22],a,q1[22]);
xor(w7[21],a,q1[21]);
xor(w7[20],a,q1[20]);
xor(w7[19],a,q1[19]);
xor(w7[18],a,q1[18]);
xor(w7[17],a,q1[17]);
xor(w7[16],a,q1[16]);
xor(w7[15],a,q1[15]);
xor(w7[14],a,q1[14]);
xor(w7[13],a,q1[13]);
xor(w7[12],a,q1[12]);
xor(w7[11],a,q1[11]);
xor(w7[10],a,q1[10]);
xor(w7[9],a,q1[9]);
xor(w7[8],a,q1[8]);
xor(w7[7],a,q1[7]);
xor(w7[6],a,q1[6]);
xor(w7[5],a,q1[5]);
xor(w7[4],a,q1[4]);
xor(w7[3],a,q1[3]);
xor(w7[2],a,q1[2]);
xor(w7[1],a,q1[1]);
//not n6(r[0],~q1[1]);
xor(w7[0],a,q1[0]);
//not n6[31:0](r,~w7[31:0]);
//not n6(r[31],~a);

halfadd ha0(q[0],w8[0],w7[0],a);
halfadd ha1(q[1],w8[1],w7[1],w8[0]);
halfadd ha2(q[2],w8[2],w7[2],w8[1]);
halfadd ha3(q[3],w8[3],w7[3],w8[2]);
halfadd ha4(q[4],w8[4],w7[4],w8[3]);
halfadd ha5(q[5],w8[5],w7[5],w8[4]);
halfadd ha6(q[6],w8[6],w7[6],w8[5]);
halfadd ha7(q[7],w8[7],w7[7],w8[6]);
halfadd ha8(q[8],w8[8],w7[8],w8[7]);
halfadd ha9(q[9],w8[9],w7[9],w8[8]);
halfadd ha10(q[10],w8[10],w7[10],w8[9]);
halfadd ha11(q[11],w8[11],w7[11],w8[10]);
halfadd ha12(q[12],w8[12],w7[12],w8[11]);
halfadd ha13(q[13],w8[13],w7[13],w8[12]);
halfadd ha14(q[14],w8[14],w7[14],w8[13]);
halfadd ha15(q[15],w8[15],w7[15],w8[14]);
halfadd ha16(q[16],w8[16],w7[16],w8[15]);
halfadd ha17(q[17],w8[17],w7[17],w8[16]);
halfadd ha18(q[18],w8[18],w7[18],w8[17]);
halfadd ha19(q[19],w8[19],w7[19],w8[18]);
halfadd ha20(q[20],w8[20],w7[20],w8[19]);
halfadd ha21(q[21],w8[21],w7[21],w8[20]);
halfadd ha22(q[22],w8[22],w7[22],w8[21]);
halfadd ha23(q[23],w8[23],w7[23],w8[22]);
halfadd ha24(q[24],w8[24],w7[24],w8[23]);
halfadd ha25(q[25],w8[25],w7[25],w8[24]);
halfadd ha26(q[26],w8[26],w7[26],w8[25]);
halfadd ha27(q[27],w8[27],w7[27],w8[26]);
halfadd ha28(q[28],w8[28],w7[28],w8[27]);
halfadd ha29(q[29],w8[29],w7[29],w8[28]);
halfadd ha30(q[30],w8[30],w7[30],w8[29]);
halfadd ha31(q[31],w8[31],w7[31],w8[30]);
//halfadd ha32(q[32],w8[32],w7[32],w8[31]);
//not n6[31:0](r,~q[31:0]);
//converting normalised form of remainder into output form//

wire b;
wire c;
not(c,m[31]);
and(b,d[31],c);
xor(w9[31],b,r1[31]);
xor(w9[30],b,r1[30]);
xor(w9[29],b,r1[29]);
xor(w9[28],b,r1[28]);
xor(w9[27],b,r1[27]);
xor(w9[26],b,r1[26]);
xor(w9[25],b,r1[25]);
xor(w9[24],b,r1[24]);
xor(w9[23],b,r1[23]);
xor(w9[22],b,r1[22]);
xor(w9[21],b,r1[21]);
xor(w9[20],b,r1[20]);
xor(w9[19],b,r1[19]);
xor(w9[18],b,r1[18]);
xor(w9[17],b,r1[17]);
xor(w9[16],b,r1[16]);
xor(w9[15],b,r1[15]);
xor(w9[14],b,r1[14]);
xor(w9[13],b,r1[13]);
xor(w9[12],b,r1[12]);
xor(w9[11],b,r1[11]);
xor(w9[10],b,r1[10]);
xor(w9[9],b,r1[9]);
xor(w9[8],b,r1[8]);
xor(w9[7],b,r1[7]);
xor(w9[6],b,r1[6]);
xor(w9[5],b,r1[5]);
xor(w9[4],b,r1[4]);
xor(w9[3],b,r1[3]);
xor(w9[2],b,r1[2]);
xor(w9[1],b,r1[1]);
xor(w9[0],b,r1[0]);
halfadd hf0(r[0],w10[0],w9[0],b);
halfadd hf1(r[1],w10[1],w9[1],w10[0]);
halfadd hf2(r[2],w10[2],w9[2],w10[1]);
halfadd hf3(r[3],w10[3],w9[3],w10[2]);
halfadd hf4(r[4],w10[4],w9[4],w10[3]);
halfadd hf5(r[5],w10[5],w9[5],w10[4]);
halfadd hf6(r[6],w10[6],w9[6],w10[5]);
halfadd hf7(r[7],w10[7],w9[7],w10[6]);
halfadd hf8(r[8],w10[8],w9[8],w10[7]);
halfadd hf9(r[9],w10[9],w9[9],w10[8]);
halfadd hf10(r[10],w10[10],w9[10],w10[9]);
halfadd hf11(r[11],w10[11],w9[11],w10[10]);
halfadd hf12(r[12],w10[12],w9[12],w10[11]);
halfadd hf13(r[13],w10[13],w9[13],w10[12]);
halfadd hf14(r[14],w10[14],w9[14],w10[13]);
halfadd hf15(r[15],w10[15],w9[15],w10[14]);
halfadd hf16(r[16],w10[16],w9[16],w10[15]);
halfadd hf17(r[17],w10[17],w9[17],w10[16]);
halfadd hf18(r[18],w10[18],w9[18],w10[17]);
halfadd hf19(r[19],w10[19],w9[19],w10[18]);
halfadd hf20(r[20],w10[20],w9[20],w10[19]);
halfadd hf21(r[21],w10[21],w9[21],w10[20]);
halfadd hf22(r[22],w10[22],w9[22],w10[21]);
halfadd hf23(r[23],w10[23],w9[23],w10[22]);
halfadd hf24(r[24],w10[24],w9[24],w10[23]);
halfadd hf25(r[25],w10[25],w9[25],w10[24]);
halfadd hf26(r[26],w10[26],w9[26],w10[25]);
halfadd hf27(r[27],w10[27],w9[27],w10[26]);
halfadd hf28(r[28],w10[28],w9[28],w10[27]);
halfadd hf29(r[29],w10[29],w9[29],w10[28]);
halfadd hf30(r[30],w10[30],w9[30],w10[29]);
halfadd hf31(r[31],w10[31],w9[31],w10[30]);

                                                    /* edhar ko change kiya */

endmodule

/*

module fulladd(sum, c_out, a, b, c_in);


output sum;
output c_out;

input a;
input b;
input c_in;

wire s1, c1, c2;


xor(s1, a, b);

xor(sum, s1, c_in);



and(c1, a, b);

and(c2, s1, c_in);


or(c_out, c2, c1);



endmodule

*/
module halfadd(sum,c_out,a,b);
output sum,c_out;
input a,b;
xor(sum,a,b);
and(c_out,a,b);
endmodule


//Define 31-bit full adder
module fulladd32bit(sum, c_out, a, b, c_in);

// I/O port declaration
output [31:0] sum;
output c_out; 
input [31:0]a;
input [31:0]b;
input c_in;

//internal nets
wire c1, c2, c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,c31;

//Instantiate four 1-bit adders
fulladd fa0(sum[0], c1, a[0], b[0], c_in);
fulladd fa1(sum[1], c2, a[1], b[1], c1);
fulladd fa2(sum[2], c3, a[2], b[2], c2);
fulladd fa3(sum[3], c4, a[3], b[3], c3);
fulladd fa4(sum[4], c5, a[4], b[4], c4);
fulladd fa5(sum[5], c6, a[5], b[5], c5);
fulladd fa6(sum[6], c7, a[6], b[6], c6);
fulladd fa7(sum[7], c8, a[7], b[7], c7);
fulladd fa8(sum[8], c9, a[8], b[8], c8);
fulladd fa9(sum[9], c10, a[9], b[9], c9);
fulladd fa10(sum[10], c11, a[10], b[10], c10);
fulladd fa11(sum[11], c12, a[11], b[11], c11);
fulladd fa12(sum[12], c13, a[12], b[12], c12);
fulladd fa13(sum[13], c14, a[13], b[13], c13);
fulladd fa14(sum[14], c15, a[14], b[14], c14);
fulladd fa15(sum[15], c16, a[15], b[15], c15);
fulladd fa16(sum[16], c17, a[16], b[16], c16);
fulladd fa17(sum[17], c18, a[17], b[17], c17);
fulladd fa18(sum[18], c19, a[18], b[18], c18);
fulladd fa19(sum[19], c20, a[19], b[19], c19);
fulladd fa20(sum[20], c21, a[20], b[20], c20);
fulladd fa21(sum[21], c22, a[21], b[21], c21);
fulladd fa22(sum[22], c23, a[22], b[22], c22);
fulladd fa23(sum[23], c24, a[23], b[23], c23);
fulladd fa24(sum[24], c25, a[24], b[24], c24);
fulladd fa25(sum[25], c26, a[25], b[25], c25);
fulladd fa26(sum[26], c27, a[26], b[26], c26);
fulladd fa27(sum[27], c28, a[27], b[27], c27);
fulladd fa28(sum[28], c29, a[28], b[28], c28);
fulladd fa29(sum[29], c30, a[29], b[29], c29);
fulladd fa30(sum[30], c31, a[30], b[30], c30);
fulladd fa31(sum[31], c_out, a[31], b[31], c31);

endmodule



module shifter(out,in,i);
output [31:0]out;
input [31:0]in;
input i;
assign out[31]=in[30];
assign out[30]=in[29];
assign out[29]=in[28];
assign out[28]=in[27];
assign out[27]=in[26];
assign out[26]=in[25];
assign out[25]=in[24];
assign out[24]=in[23];
assign out[23]=in[22];
assign out[22]=in[21];
assign out[21]=in[20];
assign out[20]=in[19];
assign out[19]=in[18];
assign out[18]=in[17];
assign out[17]=in[16];
assign out[16]=in[15];
assign out[15]=in[14];
assign out[14]=in[13];
assign out[13]=in[12];
assign out[12]=in[11];
assign out[11]=in[10];
assign out[10]=in[9];
assign out[9]=in[8];
assign out[8]=in[7];
assign out[7]=in[6];
assign out[6]=in[5];
assign out[5]=in[4];
assign out[4]=in[3];
assign out[3]=in[2];
assign out[2]=in[1];
assign out[1]=in[0];
assign out[0]=i;
endmodule


module mux(out,in1,in2,s);
output out;
input in1,in2;
input s;
wire w11,w12,w13;
not(w11,s);
and(w12,w11,in1);
and(w13,s,in2);
or(out,w12,w13);



endmodule

/*

module stimulus;
reg [31:0]m1;
reg [31:0]d1;
wire [31:0]q1;
wire [31:0]r2;

signeddivision1 sd1(q1,r2,m1,d1);
initial
begin
     $monitor($time,":\ndivisor   = %b,\ndividend  = %b\nQuotient  = %b,\nRemainder = %b", m1, d1,q1, r2);
end	 
initial
begin
         m1= 32'd14; d1=32'd15;
#5		  m1= -32'sd3; d1=32'd5;
#5       m1= 32'sd4; d1=-32'sd6;
#5       m1= -32'sd4; d1=-32'sd6;
end
endmodule	 */