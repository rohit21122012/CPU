module logic(output [31:0] LogicAnswerOne, output [31:0] LogicAnswerTwo, input [31:0] A,input [31:0] B, input S_or_U, input OpCode);

endmodule