//b12015 Rohit Patiyal 


module Logic(output [31:0] LogicAnswer, input [31:0] A,input [31:0] B, input S_or_U, input OpCode);


endmodule
