//Define 48 to 16 multiplexer
module mux48to16(out , in1 , in2 ,in3, in4 ,control,dr ,orf);

// I/O port declaration
output [31:0] out;
input [31:0] in1,in2,in3,in4;
input control,orf,dr;

//internal nets
wire control_not,fr_not;
wire [31:0] anded_out_1,anded_out_2,anded_out_3,anded_out_4;

//internal gate circuitry
not (control_not,control);
not (dr_not , dr);

and (anded_out_1[0] ,orf,dr_not, control_not , in1[0]);
and (anded_out_1[1] ,orf,dr_not, control_not , in1[1]);
and (anded_out_1[2] ,orf,dr_not, control_not , in1[2]);
and (anded_out_1[3] ,orf,dr_not, control_not , in1[3]);
and (anded_out_1[4] ,orf,dr_not, control_not , in1[4]);
and (anded_out_1[5] ,orf,dr_not, control_not , in1[5]);
and (anded_out_1[6] ,orf,dr_not, control_not , in1[6]);
and (anded_out_1[7] ,orf,dr_not, control_not , in1[7]);
and (anded_out_1[8] ,orf,dr_not, control_not , in1[8]);
and (anded_out_1[9] ,orf,dr_not, control_not , in1[9]);
and (anded_out_1[10] ,orf,dr_not, control_not , in1[10]);
and (anded_out_1[11] ,orf,dr_not, control_not , in1[11]);
and (anded_out_1[12] ,orf,dr_not, control_not , in1[12]);
and (anded_out_1[13] ,orf,dr_not, control_not , in1[13]);
and (anded_out_1[14] ,orf,dr_not, control_not , in1[14]);
and (anded_out_1[15] ,orf,dr_not, control_not , in1[15]);
and (anded_out_1[16] ,orf,dr_not, control_not , in1[16]);
and (anded_out_1[17] ,orf,dr_not, control_not , in1[17]);
and (anded_out_1[18] ,orf,dr_not, control_not , in1[18]);
and (anded_out_1[19] ,orf,dr_not, control_not , in1[19]);
and (anded_out_1[20] ,orf,dr_not, control_not , in1[20]);
and (anded_out_1[21] ,orf,dr_not, control_not , in1[21]);
and (anded_out_1[22] ,orf,dr_not, control_not , in1[22]);
and (anded_out_1[23] ,orf,dr_not, control_not , in1[23]);
and (anded_out_1[24] ,orf,dr_not, control_not , in1[24]);
and (anded_out_1[25] ,orf,dr_not, control_not , in1[25]);
and (anded_out_1[26] ,orf,dr_not, control_not , in1[26]);
and (anded_out_1[27] ,orf,dr_not, control_not , in1[27]);
and (anded_out_1[28] ,orf,dr_not, control_not , in1[28]);
and (anded_out_1[29] ,orf,dr_not, control_not , in1[29]);
and (anded_out_1[30] ,orf,dr_not, control_not , in1[30]);
and (anded_out_1[31] ,orf,dr_not, control_not , in1[31]);

and (anded_out_2[0] ,orf,dr_not, control , in2[0]);
and (anded_out_2[1] ,orf,dr_not, control , in2[1]);
and (anded_out_2[2] ,orf,dr_not, control , in2[2]);
and (anded_out_2[3] ,orf,dr_not, control , in2[3]);
and (anded_out_2[4] ,orf,dr_not, control , in2[4]);
and (anded_out_2[5] ,orf,dr_not, control , in2[5]);
and (anded_out_2[6] ,orf,dr_not, control , in2[6]);
and (anded_out_2[7] ,orf,dr_not, control , in2[7]);
and (anded_out_2[8] ,orf,dr_not, control , in2[8]);
and (anded_out_2[9] ,orf,dr_not, control , in2[9]);
and (anded_out_2[10] ,orf,dr_not, control , in2[10]);
and (anded_out_2[11] ,orf,dr_not, control , in2[11]);
and (anded_out_2[12] ,orf,dr_not, control , in2[12]);
and (anded_out_2[13] ,orf,dr_not, control , in2[13]);
and (anded_out_2[14] ,orf,dr_not, control , in2[14]);
and (anded_out_2[15] ,orf,dr_not, control , in2[15]);
and (anded_out_2[16] ,orf,dr_not, control , in2[16]);
and (anded_out_2[17] ,orf,dr_not, control , in2[17]);
and (anded_out_2[18] ,orf,dr_not, control , in2[18]);
and (anded_out_2[19] ,orf,dr_not, control , in2[19]);
and (anded_out_2[20] ,orf,dr_not, control , in2[20]);
and (anded_out_2[21] ,orf,dr_not, control , in2[21]);
and (anded_out_2[22] ,orf,dr_not, control , in2[22]);
and (anded_out_2[23] ,orf,dr_not, control , in2[23]);
and (anded_out_2[24] ,orf,dr_not, control , in2[24]);
and (anded_out_2[25] ,orf,dr_not, control , in2[25]);
and (anded_out_2[26] ,orf,dr_not, control , in2[26]);
and (anded_out_2[27] ,orf,dr_not, control , in2[27]);
and (anded_out_2[28] ,orf,dr_not, control , in2[28]);
and (anded_out_2[29] ,orf,dr_not, control , in2[29]);
and (anded_out_2[30] ,orf,dr_not, control , in2[30]);
and (anded_out_2[31] ,orf,dr_not, control , in2[31]);

and (anded_out_3[0] ,orf,dr, control_not , in3[0]);
and (anded_out_3[1] ,orf,dr, control_not , in3[1]);
and (anded_out_3[2] ,orf,dr, control_not , in3[2]);
and (anded_out_3[3] ,orf,dr, control_not , in3[3]);
and (anded_out_3[4] ,orf,dr, control_not , in3[4]);
and (anded_out_3[5] ,orf,dr, control_not , in3[5]);
and (anded_out_3[6] ,orf,dr, control_not , in3[6]);
and (anded_out_3[7] ,orf,dr, control_not , in3[7]);
and (anded_out_3[8] ,orf,dr, control_not , in3[8]);
and (anded_out_3[9] ,orf,dr, control_not , in3[9]);
and (anded_out_3[10] ,orf,dr, control_not , in3[10]);
and (anded_out_3[11] ,orf,dr, control_not , in3[11]);
and (anded_out_3[12] ,orf,dr, control_not , in3[12]);
and (anded_out_3[13] ,orf,dr, control_not , in3[13]);
and (anded_out_3[14] ,orf,dr, control_not , in3[14]);
and (anded_out_3[15] ,orf,dr, control_not , in3[15]);
and (anded_out_3[16] ,orf,dr, control_not , in3[16]);
and (anded_out_3[17] ,orf,dr, control_not , in3[17]);
and (anded_out_3[18] ,orf,dr, control_not , in3[18]);
and (anded_out_3[19] ,orf,dr, control_not , in3[19]);
and (anded_out_3[20] ,orf,dr, control_not , in3[20]);
and (anded_out_3[21] ,orf,dr, control_not , in3[21]);
and (anded_out_3[22] ,orf,dr, control_not , in3[22]);
and (anded_out_3[23] ,orf,dr, control_not , in3[23]);
and (anded_out_3[24] ,orf,dr, control_not , in3[24]);
and (anded_out_3[25] ,orf,dr, control_not , in3[25]);
and (anded_out_3[26] ,orf,dr, control_not , in3[26]);
and (anded_out_3[27] ,orf,dr, control_not , in3[27]);
and (anded_out_3[28] ,orf,dr, control_not , in3[28]);
and (anded_out_3[29] ,orf,dr, control_not , in3[29]);
and (anded_out_3[30] ,orf,dr, control_not , in3[30]);
and (anded_out_3[31] ,orf,dr, control_not , in3[31]);

and (anded_out_4[0] ,orf,dr, control , in4[0]);
and (anded_out_4[1] ,orf,dr, control , in4[1]);
and (anded_out_4[2] ,orf,dr, control , in4[2]);
and (anded_out_4[3] ,orf,dr, control , in4[3]);
and (anded_out_4[4] ,orf,dr, control , in4[4]);
and (anded_out_4[5] ,orf,dr, control , in4[5]);
and (anded_out_4[6] ,orf,dr, control , in4[6]);
and (anded_out_4[7] ,orf,dr, control , in4[7]);
and (anded_out_4[8] ,orf,dr, control , in4[8]);
and (anded_out_4[9] ,orf,dr, control , in4[9]);
and (anded_out_4[10] ,orf,dr, control , in4[10]);
and (anded_out_4[11] ,orf,dr, control , in4[11]);
and (anded_out_4[12] ,orf,dr, control , in4[12]);
and (anded_out_4[13] ,orf,dr, control , in4[13]);
and (anded_out_4[14] ,orf,dr, control , in4[14]);
and (anded_out_4[15] ,orf,dr, control , in4[15]);
and (anded_out_4[16] ,orf,dr, control , in4[16]);
and (anded_out_4[17] ,orf,dr, control , in4[17]);
and (anded_out_4[18] ,orf,dr, control , in4[18]);
and (anded_out_4[19] ,orf,dr, control , in4[19]);
and (anded_out_4[20] ,orf,dr, control , in4[20]);
and (anded_out_4[21] ,orf,dr, control , in4[21]);
and (anded_out_4[22] ,orf,dr, control , in4[22]);
and (anded_out_4[23] ,orf,dr, control , in4[23]);
and (anded_out_4[24] ,orf,dr, control , in4[24]);
and (anded_out_4[25] ,orf,dr, control , in4[25]);
and (anded_out_4[26] ,orf,dr, control , in4[26]);
and (anded_out_4[27] ,orf,dr, control , in4[27]);
and (anded_out_4[28] ,orf,dr, control , in4[28]);
and (anded_out_4[29] ,orf,dr, control , in4[29]);
and (anded_out_4[30] ,orf,dr, control , in4[30]);
and (anded_out_4[31] ,orf,dr, control , in4[31]);

or (out[0] , anded_out_1[0] , anded_out_2[0],anded_out_3[0],anded_out_4[0]);
or (out[1] , anded_out_1[1] , anded_out_2[1],anded_out_3[1],anded_out_4[1]);
or (out[2] , anded_out_1[2] , anded_out_2[2],anded_out_3[2],anded_out_4[2]);
or (out[3] , anded_out_1[3] , anded_out_2[3],anded_out_3[3],anded_out_4[3]);
or (out[4] , anded_out_1[4] , anded_out_2[4],anded_out_3[4],anded_out_4[4]);
or (out[5] , anded_out_1[5] , anded_out_2[5],anded_out_3[5],anded_out_4[5]);
or (out[6] , anded_out_1[6] , anded_out_2[6],anded_out_3[6],anded_out_4[6]);
or (out[7] , anded_out_1[7] , anded_out_2[7],anded_out_3[7],anded_out_4[7]);
or (out[8] , anded_out_1[8] , anded_out_2[8],anded_out_3[8],anded_out_4[8]);
or (out[9] , anded_out_1[9] , anded_out_2[9],anded_out_3[9],anded_out_4[9]);
or (out[10] , anded_out_1[10] , anded_out_2[10],anded_out_3[10],anded_out_4[10]);
or (out[11] , anded_out_1[11] , anded_out_2[11],anded_out_3[11],anded_out_4[11]);
or (out[12] , anded_out_1[12] , anded_out_2[12],anded_out_3[12],anded_out_4[12]);
or (out[13] , anded_out_1[13] , anded_out_2[13],anded_out_3[13],anded_out_4[13]);
or (out[14] , anded_out_1[14] , anded_out_2[14],anded_out_3[14],anded_out_4[14]);
or (out[15] , anded_out_1[15] , anded_out_2[15],anded_out_3[15],anded_out_4[15]);
or (out[16] , anded_out_1[16] , anded_out_2[16],anded_out_3[16],anded_out_4[16]);
or (out[17] , anded_out_1[17] , anded_out_2[17],anded_out_3[17],anded_out_4[17]);
or (out[18] , anded_out_1[18] , anded_out_2[18],anded_out_3[18],anded_out_4[18]);
or (out[19] , anded_out_1[19] , anded_out_2[19],anded_out_3[19],anded_out_4[19]);
or (out[20] , anded_out_1[20] , anded_out_2[20],anded_out_3[20],anded_out_4[20]);
or (out[21] , anded_out_1[21] , anded_out_2[21],anded_out_3[21],anded_out_4[21]);
or (out[22] , anded_out_1[22] , anded_out_2[22],anded_out_3[22],anded_out_4[22]);
or (out[23] , anded_out_1[23] , anded_out_2[23],anded_out_3[23],anded_out_4[23]);
or (out[24] , anded_out_1[24] , anded_out_2[24],anded_out_3[24],anded_out_4[24]);
or (out[25] , anded_out_1[25] , anded_out_2[25],anded_out_3[25],anded_out_4[25]);
or (out[26] , anded_out_1[26] , anded_out_2[26],anded_out_3[26],anded_out_4[26]);
or (out[27] , anded_out_1[27] , anded_out_2[27],anded_out_3[27],anded_out_4[27]);
or (out[28] , anded_out_1[28] , anded_out_2[28],anded_out_3[28],anded_out_4[28]);
or (out[29] , anded_out_1[29] , anded_out_2[29],anded_out_3[29],anded_out_4[29]);
or (out[30] , anded_out_1[30] , anded_out_2[30],anded_out_3[30],anded_out_4[30]);
or (out[31] , anded_out_1[31] , anded_out_2[31],anded_out_3[31],anded_out_4[31]);


endmodule